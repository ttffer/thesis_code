module layer0_cnn_121_25x64x10
(
    input clk,
    input rst,
    input [304-1:0] layer_in,
    input valid,
    output  reg ready,
    output [27*64-1:0] layer_out
);
parameter DATA_WIDTH = 27;
parameter INPUT_DATA_CNT   =   16;
reg    signed [DATA_WIDTH-1:0]  in_buffer[0:INPUT_DATA_CNT-1];
genvar j;
generate
for(j=0;j<INPUT_DATA_CNT;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=layer_in[j*19+18:j*19+0];
                    end
            end
    end
endgenerate
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=$signed(in_buffer[0]*(0));$signed(in_buffer[1]*(28));$signed(in_buffer[2]*(16));$signed(in_buffer[3]*(-32));$signed(in_buffer[4]*(4));$signed(in_buffer[5]*(-30));$signed(in_buffer[6]*(-14));$signed(in_buffer[7]*(-23));$signed(in_buffer[8]*(-10));$signed(in_buffer[9]*(7));$signed(in_buffer[10]*(-21));$signed(in_buffer[11]*(-18));$signed(in_buffer[12]*(8));$signed(in_buffer[13]*(-11));$signed(in_buffer[14]*(13));$signed(in_buffer[15]*(-27));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=$signed(in_buffer[0]*(2));$signed(in_buffer[1]*(-17));$signed(in_buffer[2]*(34));$signed(in_buffer[3]*(8));$signed(in_buffer[4]*(-13));$signed(in_buffer[5]*(-2));$signed(in_buffer[6]*(3));$signed(in_buffer[7]*(22));$signed(in_buffer[8]*(47));$signed(in_buffer[9]*(65));$signed(in_buffer[10]*(-62));$signed(in_buffer[11]*(2));$signed(in_buffer[12]*(40));$signed(in_buffer[13]*(20));$signed(in_buffer[14]*(16));$signed(in_buffer[15]*(-15));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=$signed(in_buffer[0]*(-36));$signed(in_buffer[1]*(50));$signed(in_buffer[2]*(78));$signed(in_buffer[3]*(15));$signed(in_buffer[4]*(34));$signed(in_buffer[5]*(14));$signed(in_buffer[6]*(13));$signed(in_buffer[7]*(-13));$signed(in_buffer[8]*(-18));$signed(in_buffer[9]*(-31));$signed(in_buffer[10]*(19));$signed(in_buffer[11]*(68));$signed(in_buffer[12]*(0));$signed(in_buffer[13]*(68));$signed(in_buffer[14]*(-25));$signed(in_buffer[15]*(44));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=$signed(in_buffer[0]*(21));$signed(in_buffer[1]*(-10));$signed(in_buffer[2]*(12));$signed(in_buffer[3]*(-15));$signed(in_buffer[4]*(16));$signed(in_buffer[5]*(44));$signed(in_buffer[6]*(5));$signed(in_buffer[7]*(12));$signed(in_buffer[8]*(75));$signed(in_buffer[9]*(-39));$signed(in_buffer[10]*(-8));$signed(in_buffer[11]*(20));$signed(in_buffer[12]*(6));$signed(in_buffer[13]*(33));$signed(in_buffer[14]*(-23));$signed(in_buffer[15]*(-34));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=$signed(in_buffer[0]*(5));$signed(in_buffer[1]*(-25));$signed(in_buffer[2]*(-30));$signed(in_buffer[3]*(41));$signed(in_buffer[4]*(-1));$signed(in_buffer[5]*(-9));$signed(in_buffer[6]*(-49));$signed(in_buffer[7]*(12));$signed(in_buffer[8]*(52));$signed(in_buffer[9]*(38));$signed(in_buffer[10]*(34));$signed(in_buffer[11]*(-16));$signed(in_buffer[12]*(-28));$signed(in_buffer[13]*(45));$signed(in_buffer[14]*(4));$signed(in_buffer[15]*(-25));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=$signed(in_buffer[0]*(-3));$signed(in_buffer[1]*(2));$signed(in_buffer[2]*(-19));$signed(in_buffer[3]*(17));$signed(in_buffer[4]*(-3));$signed(in_buffer[5]*(-13));$signed(in_buffer[6]*(-3));$signed(in_buffer[7]*(27));$signed(in_buffer[8]*(-25));$signed(in_buffer[9]*(-13));$signed(in_buffer[10]*(-19));$signed(in_buffer[11]*(-15));$signed(in_buffer[12]*(-24));$signed(in_buffer[13]*(-30));$signed(in_buffer[14]*(6));$signed(in_buffer[15]*(14));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=$signed(in_buffer[0]*(32));$signed(in_buffer[1]*(18));$signed(in_buffer[2]*(-21));$signed(in_buffer[3]*(-65));$signed(in_buffer[4]*(-36));$signed(in_buffer[5]*(-52));$signed(in_buffer[6]*(-52));$signed(in_buffer[7]*(-72));$signed(in_buffer[8]*(15));$signed(in_buffer[9]*(26));$signed(in_buffer[10]*(-20));$signed(in_buffer[11]*(34));$signed(in_buffer[12]*(4));$signed(in_buffer[13]*(50));$signed(in_buffer[14]*(53));$signed(in_buffer[15]*(52));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=$signed(in_buffer[0]*(-24));$signed(in_buffer[1]*(4));$signed(in_buffer[2]*(98));$signed(in_buffer[3]*(122));$signed(in_buffer[4]*(26));$signed(in_buffer[5]*(77));$signed(in_buffer[6]*(-52));$signed(in_buffer[7]*(-171));$signed(in_buffer[8]*(-1));$signed(in_buffer[9]*(-9));$signed(in_buffer[10]*(-11));$signed(in_buffer[11]*(76));$signed(in_buffer[12]*(-58));$signed(in_buffer[13]*(-2));$signed(in_buffer[14]*(-9));$signed(in_buffer[15]*(38));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=$signed(in_buffer[0]*(41));$signed(in_buffer[1]*(43));$signed(in_buffer[2]*(9));$signed(in_buffer[3]*(58));$signed(in_buffer[4]*(-34));$signed(in_buffer[5]*(-58));$signed(in_buffer[6]*(-45));$signed(in_buffer[7]*(-48));$signed(in_buffer[8]*(47));$signed(in_buffer[9]*(69));$signed(in_buffer[10]*(68));$signed(in_buffer[11]*(-26));$signed(in_buffer[12]*(32));$signed(in_buffer[13]*(-79));$signed(in_buffer[14]*(48));$signed(in_buffer[15]*(22));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=$signed(in_buffer[0]*(31));$signed(in_buffer[1]*(-55));$signed(in_buffer[2]*(-65));$signed(in_buffer[3]*(-12));$signed(in_buffer[4]*(-12));$signed(in_buffer[5]*(8));$signed(in_buffer[6]*(-61));$signed(in_buffer[7]*(-72));$signed(in_buffer[8]*(49));$signed(in_buffer[9]*(-17));$signed(in_buffer[10]*(72));$signed(in_buffer[11]*(-4));$signed(in_buffer[12]*(-48));$signed(in_buffer[13]*(19));$signed(in_buffer[14]*(38));$signed(in_buffer[15]*(-24));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight10;
assign in_buffer_weight10=$signed(in_buffer[0]*(6));$signed(in_buffer[1]*(-31));$signed(in_buffer[2]*(19));$signed(in_buffer[3]*(2));$signed(in_buffer[4]*(4));$signed(in_buffer[5]*(-14));$signed(in_buffer[6]*(-51));$signed(in_buffer[7]*(-4));$signed(in_buffer[8]*(57));$signed(in_buffer[9]*(13));$signed(in_buffer[10]*(57));$signed(in_buffer[11]*(18));$signed(in_buffer[12]*(-27));$signed(in_buffer[13]*(43));$signed(in_buffer[14]*(8));$signed(in_buffer[15]*(-41));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight11;
assign in_buffer_weight11=$signed(in_buffer[0]*(-13));$signed(in_buffer[1]*(-7));$signed(in_buffer[2]*(89));$signed(in_buffer[3]*(1));$signed(in_buffer[4]*(37));$signed(in_buffer[5]*(-41));$signed(in_buffer[6]*(22));$signed(in_buffer[7]*(74));$signed(in_buffer[8]*(-9));$signed(in_buffer[9]*(-49));$signed(in_buffer[10]*(-47));$signed(in_buffer[11]*(6));$signed(in_buffer[12]*(51));$signed(in_buffer[13]*(-22));$signed(in_buffer[14]*(-16));$signed(in_buffer[15]*(49));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight12;
assign in_buffer_weight12=$signed(in_buffer[0]*(-103));$signed(in_buffer[1]*(-3));$signed(in_buffer[2]*(18));$signed(in_buffer[3]*(71));$signed(in_buffer[4]*(-124));$signed(in_buffer[5]*(75));$signed(in_buffer[6]*(18));$signed(in_buffer[7]*(-86));$signed(in_buffer[8]*(-15));$signed(in_buffer[9]*(16));$signed(in_buffer[10]*(-19));$signed(in_buffer[11]*(-66));$signed(in_buffer[12]*(9));$signed(in_buffer[13]*(-50));$signed(in_buffer[14]*(53));$signed(in_buffer[15]*(64));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight13;
assign in_buffer_weight13=$signed(in_buffer[0]*(41));$signed(in_buffer[1]*(16));$signed(in_buffer[2]*(-16));$signed(in_buffer[3]*(49));$signed(in_buffer[4]*(-4));$signed(in_buffer[5]*(9));$signed(in_buffer[6]*(67));$signed(in_buffer[7]*(-8));$signed(in_buffer[8]*(-34));$signed(in_buffer[9]*(42));$signed(in_buffer[10]*(-4));$signed(in_buffer[11]*(14));$signed(in_buffer[12]*(-9));$signed(in_buffer[13]*(-84));$signed(in_buffer[14]*(-34));$signed(in_buffer[15]*(50));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight14;
assign in_buffer_weight14=$signed(in_buffer[0]*(-122));$signed(in_buffer[1]*(-61));$signed(in_buffer[2]*(-35));$signed(in_buffer[3]*(77));$signed(in_buffer[4]*(-152));$signed(in_buffer[5]*(-48));$signed(in_buffer[6]*(61));$signed(in_buffer[7]*(-78));$signed(in_buffer[8]*(-29));$signed(in_buffer[9]*(52));$signed(in_buffer[10]*(7));$signed(in_buffer[11]*(24));$signed(in_buffer[12]*(-43));$signed(in_buffer[13]*(34));$signed(in_buffer[14]*(-11));$signed(in_buffer[15]*(-11));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight15;
assign in_buffer_weight15=$signed(in_buffer[0]*(-1));$signed(in_buffer[1]*(9));$signed(in_buffer[2]*(21));$signed(in_buffer[3]*(-5));$signed(in_buffer[4]*(27));$signed(in_buffer[5]*(-12));$signed(in_buffer[6]*(1));$signed(in_buffer[7]*(30));$signed(in_buffer[8]*(45));$signed(in_buffer[9]*(69));$signed(in_buffer[10]*(42));$signed(in_buffer[11]*(23));$signed(in_buffer[12]*(-106));$signed(in_buffer[13]*(-74));$signed(in_buffer[14]*(1));$signed(in_buffer[15]*(-59));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight16;
assign in_buffer_weight16=$signed(in_buffer[0]*(16));$signed(in_buffer[1]*(66));$signed(in_buffer[2]*(-4));$signed(in_buffer[3]*(89));$signed(in_buffer[4]*(60));$signed(in_buffer[5]*(95));$signed(in_buffer[6]*(52));$signed(in_buffer[7]*(-12));$signed(in_buffer[8]*(9));$signed(in_buffer[9]*(4));$signed(in_buffer[10]*(-47));$signed(in_buffer[11]*(-50));$signed(in_buffer[12]*(-24));$signed(in_buffer[13]*(-18));$signed(in_buffer[14]*(-47));$signed(in_buffer[15]*(30));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight17;
assign in_buffer_weight17=$signed(in_buffer[0]*(-78));$signed(in_buffer[1]*(-74));$signed(in_buffer[2]*(-99));$signed(in_buffer[3]*(-94));$signed(in_buffer[4]*(-71));$signed(in_buffer[5]*(28));$signed(in_buffer[6]*(56));$signed(in_buffer[7]*(-15));$signed(in_buffer[8]*(4));$signed(in_buffer[9]*(-32));$signed(in_buffer[10]*(23));$signed(in_buffer[11]*(-22));$signed(in_buffer[12]*(23));$signed(in_buffer[13]*(35));$signed(in_buffer[14]*(-12));$signed(in_buffer[15]*(-17));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight18;
assign in_buffer_weight18=$signed(in_buffer[0]*(99));$signed(in_buffer[1]*(81));$signed(in_buffer[2]*(117));$signed(in_buffer[3]*(28));$signed(in_buffer[4]*(-103));$signed(in_buffer[5]*(-112));$signed(in_buffer[6]*(13));$signed(in_buffer[7]*(65));$signed(in_buffer[8]*(-12));$signed(in_buffer[9]*(-9));$signed(in_buffer[10]*(37));$signed(in_buffer[11]*(17));$signed(in_buffer[12]*(22));$signed(in_buffer[13]*(-30));$signed(in_buffer[14]*(17));$signed(in_buffer[15]*(-64));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight19;
assign in_buffer_weight19=$signed(in_buffer[0]*(-25));$signed(in_buffer[1]*(19));$signed(in_buffer[2]*(22));$signed(in_buffer[3]*(33));$signed(in_buffer[4]*(107));$signed(in_buffer[5]*(-36));$signed(in_buffer[6]*(-29));$signed(in_buffer[7]*(26));$signed(in_buffer[8]*(35));$signed(in_buffer[9]*(74));$signed(in_buffer[10]*(-2));$signed(in_buffer[11]*(-1));$signed(in_buffer[12]*(-57));$signed(in_buffer[13]*(-7));$signed(in_buffer[14]*(-40));$signed(in_buffer[15]*(17));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight20;
assign in_buffer_weight20=$signed(in_buffer[0]*(3));$signed(in_buffer[1]*(-2));$signed(in_buffer[2]*(40));$signed(in_buffer[3]*(-59));$signed(in_buffer[4]*(-28));$signed(in_buffer[5]*(21));$signed(in_buffer[6]*(-4));$signed(in_buffer[7]*(-7));$signed(in_buffer[8]*(58));$signed(in_buffer[9]*(22));$signed(in_buffer[10]*(46));$signed(in_buffer[11]*(92));$signed(in_buffer[12]*(-13));$signed(in_buffer[13]*(-45));$signed(in_buffer[14]*(-15));$signed(in_buffer[15]*(2));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight21;
assign in_buffer_weight21=$signed(in_buffer[0]*(-36));$signed(in_buffer[1]*(-15));$signed(in_buffer[2]*(-1));$signed(in_buffer[3]*(28));$signed(in_buffer[4]*(82));$signed(in_buffer[5]*(49));$signed(in_buffer[6]*(5));$signed(in_buffer[7]*(-18));$signed(in_buffer[8]*(-180));$signed(in_buffer[9]*(-76));$signed(in_buffer[10]*(36));$signed(in_buffer[11]*(-7));$signed(in_buffer[12]*(53));$signed(in_buffer[13]*(10));$signed(in_buffer[14]*(44));$signed(in_buffer[15]*(1));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight22;
assign in_buffer_weight22=$signed(in_buffer[0]*(59));$signed(in_buffer[1]*(36));$signed(in_buffer[2]*(-2));$signed(in_buffer[3]*(11));$signed(in_buffer[4]*(-23));$signed(in_buffer[5]*(-30));$signed(in_buffer[6]*(-28));$signed(in_buffer[7]*(-20));$signed(in_buffer[8]*(-47));$signed(in_buffer[9]*(21));$signed(in_buffer[10]*(5));$signed(in_buffer[11]*(-35));$signed(in_buffer[12]*(-19));$signed(in_buffer[13]*(79));$signed(in_buffer[14]*(25));$signed(in_buffer[15]*(61));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight23;
assign in_buffer_weight23=$signed(in_buffer[0]*(-100));$signed(in_buffer[1]*(-184));$signed(in_buffer[2]*(-44));$signed(in_buffer[3]*(-53));$signed(in_buffer[4]*(14));$signed(in_buffer[5]*(37));$signed(in_buffer[6]*(-19));$signed(in_buffer[7]*(34));$signed(in_buffer[8]*(83));$signed(in_buffer[9]*(38));$signed(in_buffer[10]*(7));$signed(in_buffer[11]*(21));$signed(in_buffer[12]*(-54));$signed(in_buffer[13]*(-41));$signed(in_buffer[14]*(23));$signed(in_buffer[15]*(-26));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight24;
assign in_buffer_weight24=$signed(in_buffer[0]*(68));$signed(in_buffer[1]*(105));$signed(in_buffer[2]*(49));$signed(in_buffer[3]*(-45));$signed(in_buffer[4]*(23));$signed(in_buffer[5]*(-50));$signed(in_buffer[6]*(-9));$signed(in_buffer[7]*(-1));$signed(in_buffer[8]*(-58));$signed(in_buffer[9]*(16));$signed(in_buffer[10]*(62));$signed(in_buffer[11]*(-70));$signed(in_buffer[12]*(60));$signed(in_buffer[13]*(-36));$signed(in_buffer[14]*(-17));$signed(in_buffer[15]*(10));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight25;
assign in_buffer_weight25=$signed(in_buffer[0]*(-1));$signed(in_buffer[1]*(65));$signed(in_buffer[2]*(53));$signed(in_buffer[3]*(17));$signed(in_buffer[4]*(10));$signed(in_buffer[5]*(-70));$signed(in_buffer[6]*(65));$signed(in_buffer[7]*(12));$signed(in_buffer[8]*(-37));$signed(in_buffer[9]*(-41));$signed(in_buffer[10]*(-40));$signed(in_buffer[11]*(-25));$signed(in_buffer[12]*(-6));$signed(in_buffer[13]*(89));$signed(in_buffer[14]*(-47));$signed(in_buffer[15]*(-12));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight26;
assign in_buffer_weight26=$signed(in_buffer[0]*(17));$signed(in_buffer[1]*(-2));$signed(in_buffer[2]*(7));$signed(in_buffer[3]*(15));$signed(in_buffer[4]*(-12));$signed(in_buffer[5]*(-9));$signed(in_buffer[6]*(-4));$signed(in_buffer[7]*(18));$signed(in_buffer[8]*(-35));$signed(in_buffer[9]*(-6));$signed(in_buffer[10]*(-29));$signed(in_buffer[11]*(-3));$signed(in_buffer[12]*(0));$signed(in_buffer[13]*(-9));$signed(in_buffer[14]*(-23));$signed(in_buffer[15]*(-16));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight27;
assign in_buffer_weight27=$signed(in_buffer[0]*(-71));$signed(in_buffer[1]*(-58));$signed(in_buffer[2]*(79));$signed(in_buffer[3]*(-49));$signed(in_buffer[4]*(11));$signed(in_buffer[5]*(45));$signed(in_buffer[6]*(62));$signed(in_buffer[7]*(43));$signed(in_buffer[8]*(-25));$signed(in_buffer[9]*(-53));$signed(in_buffer[10]*(43));$signed(in_buffer[11]*(55));$signed(in_buffer[12]*(-48));$signed(in_buffer[13]*(-14));$signed(in_buffer[14]*(-33));$signed(in_buffer[15]*(-80));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight28;
assign in_buffer_weight28=$signed(in_buffer[0]*(84));$signed(in_buffer[1]*(-11));$signed(in_buffer[2]*(-66));$signed(in_buffer[3]*(-1));$signed(in_buffer[4]*(129));$signed(in_buffer[5]*(-21));$signed(in_buffer[6]*(-41));$signed(in_buffer[7]*(52));$signed(in_buffer[8]*(-96));$signed(in_buffer[9]*(-13));$signed(in_buffer[10]*(8));$signed(in_buffer[11]*(-30));$signed(in_buffer[12]*(12));$signed(in_buffer[13]*(36));$signed(in_buffer[14]*(34));$signed(in_buffer[15]*(-14));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight29;
assign in_buffer_weight29=$signed(in_buffer[0]*(27));$signed(in_buffer[1]*(-6));$signed(in_buffer[2]*(20));$signed(in_buffer[3]*(20));$signed(in_buffer[4]*(8));$signed(in_buffer[5]*(-26));$signed(in_buffer[6]*(-38));$signed(in_buffer[7]*(40));$signed(in_buffer[8]*(-8));$signed(in_buffer[9]*(55));$signed(in_buffer[10]*(4));$signed(in_buffer[11]*(17));$signed(in_buffer[12]*(6));$signed(in_buffer[13]*(57));$signed(in_buffer[14]*(-38));$signed(in_buffer[15]*(32));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight30;
assign in_buffer_weight30=$signed(in_buffer[0]*(-19));$signed(in_buffer[1]*(-16));$signed(in_buffer[2]*(39));$signed(in_buffer[3]*(-28));$signed(in_buffer[4]*(11));$signed(in_buffer[5]*(37));$signed(in_buffer[6]*(19));$signed(in_buffer[7]*(-8));$signed(in_buffer[8]*(-1));$signed(in_buffer[9]*(-39));$signed(in_buffer[10]*(-13));$signed(in_buffer[11]*(55));$signed(in_buffer[12]*(0));$signed(in_buffer[13]*(59));$signed(in_buffer[14]*(-2));$signed(in_buffer[15]*(11));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight31;
assign in_buffer_weight31=$signed(in_buffer[0]*(31));$signed(in_buffer[1]*(-20));$signed(in_buffer[2]*(-58));$signed(in_buffer[3]*(-4));$signed(in_buffer[4]*(26));$signed(in_buffer[5]*(53));$signed(in_buffer[6]*(23));$signed(in_buffer[7]*(72));$signed(in_buffer[8]*(78));$signed(in_buffer[9]*(26));$signed(in_buffer[10]*(-78));$signed(in_buffer[11]*(-22));$signed(in_buffer[12]*(-25));$signed(in_buffer[13]*(-56));$signed(in_buffer[14]*(-46));$signed(in_buffer[15]*(-14));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight32;
assign in_buffer_weight32=$signed(in_buffer[0]*(-12));$signed(in_buffer[1]*(-25));$signed(in_buffer[2]*(87));$signed(in_buffer[3]*(2));$signed(in_buffer[4]*(73));$signed(in_buffer[5]*(25));$signed(in_buffer[6]*(-73));$signed(in_buffer[7]*(17));$signed(in_buffer[8]*(18));$signed(in_buffer[9]*(43));$signed(in_buffer[10]*(13));$signed(in_buffer[11]*(-4));$signed(in_buffer[12]*(-13));$signed(in_buffer[13]*(43));$signed(in_buffer[14]*(-18));$signed(in_buffer[15]*(4));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight33;
assign in_buffer_weight33=$signed(in_buffer[0]*(45));$signed(in_buffer[1]*(-6));$signed(in_buffer[2]*(8));$signed(in_buffer[3]*(-2));$signed(in_buffer[4]*(-55));$signed(in_buffer[5]*(18));$signed(in_buffer[6]*(16));$signed(in_buffer[7]*(-1));$signed(in_buffer[8]*(84));$signed(in_buffer[9]*(22));$signed(in_buffer[10]*(-6));$signed(in_buffer[11]*(109));$signed(in_buffer[12]*(-41));$signed(in_buffer[13]*(-12));$signed(in_buffer[14]*(31));$signed(in_buffer[15]*(3));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight34;
assign in_buffer_weight34=$signed(in_buffer[0]*(61));$signed(in_buffer[1]*(32));$signed(in_buffer[2]*(0));$signed(in_buffer[3]*(24));$signed(in_buffer[4]*(25));$signed(in_buffer[5]*(67));$signed(in_buffer[6]*(57));$signed(in_buffer[7]*(67));$signed(in_buffer[8]*(30));$signed(in_buffer[9]*(-47));$signed(in_buffer[10]*(-48));$signed(in_buffer[11]*(-43));$signed(in_buffer[12]*(-62));$signed(in_buffer[13]*(34));$signed(in_buffer[14]*(-46));$signed(in_buffer[15]*(-71));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight35;
assign in_buffer_weight35=$signed(in_buffer[0]*(15));$signed(in_buffer[1]*(29));$signed(in_buffer[2]*(28));$signed(in_buffer[3]*(52));$signed(in_buffer[4]*(46));$signed(in_buffer[5]*(-32));$signed(in_buffer[6]*(-26));$signed(in_buffer[7]*(-42));$signed(in_buffer[8]*(40));$signed(in_buffer[9]*(28));$signed(in_buffer[10]*(79));$signed(in_buffer[11]*(49));$signed(in_buffer[12]*(-35));$signed(in_buffer[13]*(-74));$signed(in_buffer[14]*(31));$signed(in_buffer[15]*(1));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight36;
assign in_buffer_weight36=$signed(in_buffer[0]*(10));$signed(in_buffer[1]*(29));$signed(in_buffer[2]*(-1));$signed(in_buffer[3]*(0));$signed(in_buffer[4]*(-31));$signed(in_buffer[5]*(-8));$signed(in_buffer[6]*(29));$signed(in_buffer[7]*(2));$signed(in_buffer[8]*(-17));$signed(in_buffer[9]*(1));$signed(in_buffer[10]*(-14));$signed(in_buffer[11]*(-32));$signed(in_buffer[12]*(1));$signed(in_buffer[13]*(-24));$signed(in_buffer[14]*(-33));$signed(in_buffer[15]*(-14));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight37;
assign in_buffer_weight37=$signed(in_buffer[0]*(45));$signed(in_buffer[1]*(49));$signed(in_buffer[2]*(-36));$signed(in_buffer[3]*(53));$signed(in_buffer[4]*(26));$signed(in_buffer[5]*(8));$signed(in_buffer[6]*(68));$signed(in_buffer[7]*(-16));$signed(in_buffer[8]*(-42));$signed(in_buffer[9]*(10));$signed(in_buffer[10]*(-34));$signed(in_buffer[11]*(45));$signed(in_buffer[12]*(-19));$signed(in_buffer[13]*(-53));$signed(in_buffer[14]*(-19));$signed(in_buffer[15]*(33));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight38;
assign in_buffer_weight38=$signed(in_buffer[0]*(32));$signed(in_buffer[1]*(-22));$signed(in_buffer[2]*(0));$signed(in_buffer[3]*(-6));$signed(in_buffer[4]*(-13));$signed(in_buffer[5]*(-12));$signed(in_buffer[6]*(-6));$signed(in_buffer[7]*(9));$signed(in_buffer[8]*(-28));$signed(in_buffer[9]*(-24));$signed(in_buffer[10]*(-16));$signed(in_buffer[11]*(24));$signed(in_buffer[12]*(-16));$signed(in_buffer[13]*(-27));$signed(in_buffer[14]*(22));$signed(in_buffer[15]*(4));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight39;
assign in_buffer_weight39=$signed(in_buffer[0]*(55));$signed(in_buffer[1]*(-14));$signed(in_buffer[2]*(-17));$signed(in_buffer[3]*(50));$signed(in_buffer[4]*(-14));$signed(in_buffer[5]*(1));$signed(in_buffer[6]*(-56));$signed(in_buffer[7]*(25));$signed(in_buffer[8]*(76));$signed(in_buffer[9]*(4));$signed(in_buffer[10]*(-1));$signed(in_buffer[11]*(29));$signed(in_buffer[12]*(17));$signed(in_buffer[13]*(31));$signed(in_buffer[14]*(23));$signed(in_buffer[15]*(3));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight40;
assign in_buffer_weight40=$signed(in_buffer[0]*(-15));$signed(in_buffer[1]*(8));$signed(in_buffer[2]*(9));$signed(in_buffer[3]*(-13));$signed(in_buffer[4]*(20));$signed(in_buffer[5]*(63));$signed(in_buffer[6]*(52));$signed(in_buffer[7]*(30));$signed(in_buffer[8]*(-55));$signed(in_buffer[9]*(0));$signed(in_buffer[10]*(8));$signed(in_buffer[11]*(34));$signed(in_buffer[12]*(-12));$signed(in_buffer[13]*(-11));$signed(in_buffer[14]*(-46));$signed(in_buffer[15]*(-2));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight41;
assign in_buffer_weight41=$signed(in_buffer[0]*(34));$signed(in_buffer[1]*(34));$signed(in_buffer[2]*(-5));$signed(in_buffer[3]*(-16));$signed(in_buffer[4]*(-6));$signed(in_buffer[5]*(-26));$signed(in_buffer[6]*(86));$signed(in_buffer[7]*(0));$signed(in_buffer[8]*(-9));$signed(in_buffer[9]*(-7));$signed(in_buffer[10]*(-22));$signed(in_buffer[11]*(21));$signed(in_buffer[12]*(29));$signed(in_buffer[13]*(-45));$signed(in_buffer[14]*(16));$signed(in_buffer[15]*(88));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight42;
assign in_buffer_weight42=$signed(in_buffer[0]*(-1));$signed(in_buffer[1]*(22));$signed(in_buffer[2]*(27));$signed(in_buffer[3]*(-11));$signed(in_buffer[4]*(3));$signed(in_buffer[5]*(16));$signed(in_buffer[6]*(39));$signed(in_buffer[7]*(38));$signed(in_buffer[8]*(-50));$signed(in_buffer[9]*(42));$signed(in_buffer[10]*(-41));$signed(in_buffer[11]*(11));$signed(in_buffer[12]*(73));$signed(in_buffer[13]*(-30));$signed(in_buffer[14]*(11));$signed(in_buffer[15]*(1));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight43;
assign in_buffer_weight43=$signed(in_buffer[0]*(-18));$signed(in_buffer[1]*(35));$signed(in_buffer[2]*(1));$signed(in_buffer[3]*(-84));$signed(in_buffer[4]*(-19));$signed(in_buffer[5]*(21));$signed(in_buffer[6]*(43));$signed(in_buffer[7]*(-95));$signed(in_buffer[8]*(6));$signed(in_buffer[9]*(-47));$signed(in_buffer[10]*(64));$signed(in_buffer[11]*(-25));$signed(in_buffer[12]*(-104));$signed(in_buffer[13]*(61));$signed(in_buffer[14]*(8));$signed(in_buffer[15]*(-33));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight44;
assign in_buffer_weight44=$signed(in_buffer[0]*(19));$signed(in_buffer[1]*(-9));$signed(in_buffer[2]*(61));$signed(in_buffer[3]*(-11));$signed(in_buffer[4]*(7));$signed(in_buffer[5]*(29));$signed(in_buffer[6]*(20));$signed(in_buffer[7]*(12));$signed(in_buffer[8]*(31));$signed(in_buffer[9]*(-12));$signed(in_buffer[10]*(-119));$signed(in_buffer[11]*(-21));$signed(in_buffer[12]*(67));$signed(in_buffer[13]*(-20));$signed(in_buffer[14]*(12));$signed(in_buffer[15]*(35));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight45;
assign in_buffer_weight45=$signed(in_buffer[0]*(-84));$signed(in_buffer[1]*(37));$signed(in_buffer[2]*(-17));$signed(in_buffer[3]*(36));$signed(in_buffer[4]*(-10));$signed(in_buffer[5]*(7));$signed(in_buffer[6]*(68));$signed(in_buffer[7]*(62));$signed(in_buffer[8]*(-67));$signed(in_buffer[9]*(-3));$signed(in_buffer[10]*(48));$signed(in_buffer[11]*(-39));$signed(in_buffer[12]*(25));$signed(in_buffer[13]*(16));$signed(in_buffer[14]*(-36));$signed(in_buffer[15]*(-106));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight46;
assign in_buffer_weight46=$signed(in_buffer[0]*(-75));$signed(in_buffer[1]*(10));$signed(in_buffer[2]*(31));$signed(in_buffer[3]*(29));$signed(in_buffer[4]*(-17));$signed(in_buffer[5]*(36));$signed(in_buffer[6]*(23));$signed(in_buffer[7]*(53));$signed(in_buffer[8]*(-5));$signed(in_buffer[9]*(58));$signed(in_buffer[10]*(-2));$signed(in_buffer[11]*(-57));$signed(in_buffer[12]*(60));$signed(in_buffer[13]*(-14));$signed(in_buffer[14]*(-35));$signed(in_buffer[15]*(25));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight47;
assign in_buffer_weight47=$signed(in_buffer[0]*(-1));$signed(in_buffer[1]*(-99));$signed(in_buffer[2]*(-38));$signed(in_buffer[3]*(-16));$signed(in_buffer[4]*(-128));$signed(in_buffer[5]*(-66));$signed(in_buffer[6]*(-66));$signed(in_buffer[7]*(-59));$signed(in_buffer[8]*(49));$signed(in_buffer[9]*(33));$signed(in_buffer[10]*(10));$signed(in_buffer[11]*(-12));$signed(in_buffer[12]*(49));$signed(in_buffer[13]*(32));$signed(in_buffer[14]*(73));$signed(in_buffer[15]*(79));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight48;
assign in_buffer_weight48=$signed(in_buffer[0]*(60));$signed(in_buffer[1]*(26));$signed(in_buffer[2]*(-41));$signed(in_buffer[3]*(45));$signed(in_buffer[4]*(-13));$signed(in_buffer[5]*(-45));$signed(in_buffer[6]*(-13));$signed(in_buffer[7]*(16));$signed(in_buffer[8]*(-24));$signed(in_buffer[9]*(85));$signed(in_buffer[10]*(78));$signed(in_buffer[11]*(-2));$signed(in_buffer[12]*(-106));$signed(in_buffer[13]*(-43));$signed(in_buffer[14]*(17));$signed(in_buffer[15]*(-130));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight49;
assign in_buffer_weight49=$signed(in_buffer[0]*(-125));$signed(in_buffer[1]*(-124));$signed(in_buffer[2]*(114));$signed(in_buffer[3]*(19));$signed(in_buffer[4]*(-29));$signed(in_buffer[5]*(-55));$signed(in_buffer[6]*(33));$signed(in_buffer[7]*(7));$signed(in_buffer[8]*(60));$signed(in_buffer[9]*(-30));$signed(in_buffer[10]*(8));$signed(in_buffer[11]*(32));$signed(in_buffer[12]*(30));$signed(in_buffer[13]*(29));$signed(in_buffer[14]*(4));$signed(in_buffer[15]*(-15));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight50;
assign in_buffer_weight50=$signed(in_buffer[0]*(7));$signed(in_buffer[1]*(-33));$signed(in_buffer[2]*(-12));$signed(in_buffer[3]*(-95));$signed(in_buffer[4]*(9));$signed(in_buffer[5]*(-70));$signed(in_buffer[6]*(8));$signed(in_buffer[7]*(-43));$signed(in_buffer[8]*(63));$signed(in_buffer[9]*(10));$signed(in_buffer[10]*(67));$signed(in_buffer[11]*(-31));$signed(in_buffer[12]*(38));$signed(in_buffer[13]*(22));$signed(in_buffer[14]*(-4));$signed(in_buffer[15]*(-97));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight51;
assign in_buffer_weight51=$signed(in_buffer[0]*(13));$signed(in_buffer[1]*(28));$signed(in_buffer[2]*(-18));$signed(in_buffer[3]*(29));$signed(in_buffer[4]*(57));$signed(in_buffer[5]*(-26));$signed(in_buffer[6]*(10));$signed(in_buffer[7]*(-5));$signed(in_buffer[8]*(-69));$signed(in_buffer[9]*(58));$signed(in_buffer[10]*(54));$signed(in_buffer[11]*(-56));$signed(in_buffer[12]*(-9));$signed(in_buffer[13]*(46));$signed(in_buffer[14]*(-18));$signed(in_buffer[15]*(31));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight52;
assign in_buffer_weight52=$signed(in_buffer[0]*(46));$signed(in_buffer[1]*(42));$signed(in_buffer[2]*(-26));$signed(in_buffer[3]*(-28));$signed(in_buffer[4]*(-5));$signed(in_buffer[5]*(2));$signed(in_buffer[6]*(25));$signed(in_buffer[7]*(66));$signed(in_buffer[8]*(-10));$signed(in_buffer[9]*(27));$signed(in_buffer[10]*(-59));$signed(in_buffer[11]*(7));$signed(in_buffer[12]*(12));$signed(in_buffer[13]*(6));$signed(in_buffer[14]*(-59));$signed(in_buffer[15]*(52));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight53;
assign in_buffer_weight53=$signed(in_buffer[0]*(11));$signed(in_buffer[1]*(-20));$signed(in_buffer[2]*(-26));$signed(in_buffer[3]*(-20));$signed(in_buffer[4]*(25));$signed(in_buffer[5]*(-18));$signed(in_buffer[6]*(-9));$signed(in_buffer[7]*(-25));$signed(in_buffer[8]*(16));$signed(in_buffer[9]*(-22));$signed(in_buffer[10]*(-28));$signed(in_buffer[11]*(-19));$signed(in_buffer[12]*(-20));$signed(in_buffer[13]*(4));$signed(in_buffer[14]*(8));$signed(in_buffer[15]*(-15));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight54;
assign in_buffer_weight54=$signed(in_buffer[0]*(-2));$signed(in_buffer[1]*(-127));$signed(in_buffer[2]*(-178));$signed(in_buffer[3]*(-138));$signed(in_buffer[4]*(-10));$signed(in_buffer[5]*(9));$signed(in_buffer[6]*(37));$signed(in_buffer[7]*(30));$signed(in_buffer[8]*(30));$signed(in_buffer[9]*(-26));$signed(in_buffer[10]*(-19));$signed(in_buffer[11]*(12));$signed(in_buffer[12]*(13));$signed(in_buffer[13]*(-28));$signed(in_buffer[14]*(16));$signed(in_buffer[15]*(36));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight55;
assign in_buffer_weight55=$signed(in_buffer[0]*(-65));$signed(in_buffer[1]*(-27));$signed(in_buffer[2]*(75));$signed(in_buffer[3]*(78));$signed(in_buffer[4]*(-12));$signed(in_buffer[5]*(29));$signed(in_buffer[6]*(-3));$signed(in_buffer[7]*(52));$signed(in_buffer[8]*(48));$signed(in_buffer[9]*(57));$signed(in_buffer[10]*(-27));$signed(in_buffer[11]*(-19));$signed(in_buffer[12]*(-20));$signed(in_buffer[13]*(-32));$signed(in_buffer[14]*(-29));$signed(in_buffer[15]*(15));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight56;
assign in_buffer_weight56=$signed(in_buffer[0]*(-38));$signed(in_buffer[1]*(26));$signed(in_buffer[2]*(91));$signed(in_buffer[3]*(-31));$signed(in_buffer[4]*(52));$signed(in_buffer[5]*(20));$signed(in_buffer[6]*(9));$signed(in_buffer[7]*(-40));$signed(in_buffer[8]*(17));$signed(in_buffer[9]*(-9));$signed(in_buffer[10]*(-76));$signed(in_buffer[11]*(15));$signed(in_buffer[12]*(23));$signed(in_buffer[13]*(43));$signed(in_buffer[14]*(-31));$signed(in_buffer[15]*(44));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight57;
assign in_buffer_weight57=$signed(in_buffer[0]*(-8));$signed(in_buffer[1]*(7));$signed(in_buffer[2]*(4));$signed(in_buffer[3]*(24));$signed(in_buffer[4]*(-12));$signed(in_buffer[5]*(15));$signed(in_buffer[6]*(-17));$signed(in_buffer[7]*(-3));$signed(in_buffer[8]*(15));$signed(in_buffer[9]*(-17));$signed(in_buffer[10]*(-24));$signed(in_buffer[11]*(-32));$signed(in_buffer[12]*(-13));$signed(in_buffer[13]*(-21));$signed(in_buffer[14]*(17));$signed(in_buffer[15]*(-3));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight58;
assign in_buffer_weight58=$signed(in_buffer[0]*(-30));$signed(in_buffer[1]*(6));$signed(in_buffer[2]*(-12));$signed(in_buffer[3]*(-8));$signed(in_buffer[4]*(46));$signed(in_buffer[5]*(50));$signed(in_buffer[6]*(-38));$signed(in_buffer[7]*(1));$signed(in_buffer[8]*(-71));$signed(in_buffer[9]*(24));$signed(in_buffer[10]*(53));$signed(in_buffer[11]*(-87));$signed(in_buffer[12]*(21));$signed(in_buffer[13]*(42));$signed(in_buffer[14]*(54));$signed(in_buffer[15]*(-61));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight59;
assign in_buffer_weight59=$signed(in_buffer[0]*(-23));$signed(in_buffer[1]*(22));$signed(in_buffer[2]*(8));$signed(in_buffer[3]*(15));$signed(in_buffer[4]*(-68));$signed(in_buffer[5]*(-11));$signed(in_buffer[6]*(9));$signed(in_buffer[7]*(-37));$signed(in_buffer[8]*(40));$signed(in_buffer[9]*(-73));$signed(in_buffer[10]*(-37));$signed(in_buffer[11]*(-29));$signed(in_buffer[12]*(65));$signed(in_buffer[13]*(55));$signed(in_buffer[14]*(54));$signed(in_buffer[15]*(72));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight60;
assign in_buffer_weight60=$signed(in_buffer[0]*(-89));$signed(in_buffer[1]*(-11));$signed(in_buffer[2]*(-91));$signed(in_buffer[3]*(-20));$signed(in_buffer[4]*(-76));$signed(in_buffer[5]*(-68));$signed(in_buffer[6]*(-7));$signed(in_buffer[7]*(34));$signed(in_buffer[8]*(-23));$signed(in_buffer[9]*(61));$signed(in_buffer[10]*(-25));$signed(in_buffer[11]*(-67));$signed(in_buffer[12]*(-17));$signed(in_buffer[13]*(64));$signed(in_buffer[14]*(12));$signed(in_buffer[15]*(-76));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight61;
assign in_buffer_weight61=$signed(in_buffer[0]*(28));$signed(in_buffer[1]*(59));$signed(in_buffer[2]*(53));$signed(in_buffer[3]*(2));$signed(in_buffer[4]*(12));$signed(in_buffer[5]*(43));$signed(in_buffer[6]*(-35));$signed(in_buffer[7]*(35));$signed(in_buffer[8]*(-115));$signed(in_buffer[9]*(49));$signed(in_buffer[10]*(7));$signed(in_buffer[11]*(-57));$signed(in_buffer[12]*(71));$signed(in_buffer[13]*(-26));$signed(in_buffer[14]*(-29));$signed(in_buffer[15]*(13));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight62;
assign in_buffer_weight62=$signed(in_buffer[0]*(-44));$signed(in_buffer[1]*(-73));$signed(in_buffer[2]*(-70));$signed(in_buffer[3]*(-22));$signed(in_buffer[4]*(98));$signed(in_buffer[5]*(78));$signed(in_buffer[6]*(58));$signed(in_buffer[7]*(-51));$signed(in_buffer[8]*(0));$signed(in_buffer[9]*(-13));$signed(in_buffer[10]*(39));$signed(in_buffer[11]*(-2));$signed(in_buffer[12]*(-52));$signed(in_buffer[13]*(-9));$signed(in_buffer[14]*(29));$signed(in_buffer[15]*(-53));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight63;
assign in_buffer_weight63=$signed(in_buffer[0]*(-63));$signed(in_buffer[1]*(-86));$signed(in_buffer[2]*(-22));$signed(in_buffer[3]*(74));$signed(in_buffer[4]*(-56));$signed(in_buffer[5]*(7));$signed(in_buffer[6]*(35));$signed(in_buffer[7]*(42));$signed(in_buffer[8]*(-64));$signed(in_buffer[9]*(59));$signed(in_buffer[10]*(58));$signed(in_buffer[11]*(-132));$signed(in_buffer[12]*(-26));$signed(in_buffer[13]*(-14));$signed(in_buffer[14]*(-10));$signed(in_buffer[15]*(-16));;
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
wire signed [DATA_WIDTH-1:0]   weight_bias10;
wire signed [DATA_WIDTH-1:0]   weight_bias11;
wire signed [DATA_WIDTH-1:0]   weight_bias12;
wire signed [DATA_WIDTH-1:0]   weight_bias13;
wire signed [DATA_WIDTH-1:0]   weight_bias14;
wire signed [DATA_WIDTH-1:0]   weight_bias15;
wire signed [DATA_WIDTH-1:0]   weight_bias16;
wire signed [DATA_WIDTH-1:0]   weight_bias17;
wire signed [DATA_WIDTH-1:0]   weight_bias18;
wire signed [DATA_WIDTH-1:0]   weight_bias19;
wire signed [DATA_WIDTH-1:0]   weight_bias20;
wire signed [DATA_WIDTH-1:0]   weight_bias21;
wire signed [DATA_WIDTH-1:0]   weight_bias22;
wire signed [DATA_WIDTH-1:0]   weight_bias23;
wire signed [DATA_WIDTH-1:0]   weight_bias24;
wire signed [DATA_WIDTH-1:0]   weight_bias25;
wire signed [DATA_WIDTH-1:0]   weight_bias26;
wire signed [DATA_WIDTH-1:0]   weight_bias27;
wire signed [DATA_WIDTH-1:0]   weight_bias28;
wire signed [DATA_WIDTH-1:0]   weight_bias29;
wire signed [DATA_WIDTH-1:0]   weight_bias30;
wire signed [DATA_WIDTH-1:0]   weight_bias31;
wire signed [DATA_WIDTH-1:0]   weight_bias32;
wire signed [DATA_WIDTH-1:0]   weight_bias33;
wire signed [DATA_WIDTH-1:0]   weight_bias34;
wire signed [DATA_WIDTH-1:0]   weight_bias35;
wire signed [DATA_WIDTH-1:0]   weight_bias36;
wire signed [DATA_WIDTH-1:0]   weight_bias37;
wire signed [DATA_WIDTH-1:0]   weight_bias38;
wire signed [DATA_WIDTH-1:0]   weight_bias39;
wire signed [DATA_WIDTH-1:0]   weight_bias40;
wire signed [DATA_WIDTH-1:0]   weight_bias41;
wire signed [DATA_WIDTH-1:0]   weight_bias42;
wire signed [DATA_WIDTH-1:0]   weight_bias43;
wire signed [DATA_WIDTH-1:0]   weight_bias44;
wire signed [DATA_WIDTH-1:0]   weight_bias45;
wire signed [DATA_WIDTH-1:0]   weight_bias46;
wire signed [DATA_WIDTH-1:0]   weight_bias47;
wire signed [DATA_WIDTH-1:0]   weight_bias48;
wire signed [DATA_WIDTH-1:0]   weight_bias49;
wire signed [DATA_WIDTH-1:0]   weight_bias50;
wire signed [DATA_WIDTH-1:0]   weight_bias51;
wire signed [DATA_WIDTH-1:0]   weight_bias52;
wire signed [DATA_WIDTH-1:0]   weight_bias53;
wire signed [DATA_WIDTH-1:0]   weight_bias54;
wire signed [DATA_WIDTH-1:0]   weight_bias55;
wire signed [DATA_WIDTH-1:0]   weight_bias56;
wire signed [DATA_WIDTH-1:0]   weight_bias57;
wire signed [DATA_WIDTH-1:0]   weight_bias58;
wire signed [DATA_WIDTH-1:0]   weight_bias59;
wire signed [DATA_WIDTH-1:0]   weight_bias60;
wire signed [DATA_WIDTH-1:0]   weight_bias61;
wire signed [DATA_WIDTH-1:0]   weight_bias62;
wire signed [DATA_WIDTH-1:0]   weight_bias63;
assign weight_bias0=in_buffer_weight0+(-19);
assign weight_bias1=in_buffer_weight1+(13);
assign weight_bias2=in_buffer_weight2+(-67);
assign weight_bias3=in_buffer_weight3+(72);
assign weight_bias4=in_buffer_weight4+(66);
assign weight_bias5=in_buffer_weight5+(-2);
assign weight_bias6=in_buffer_weight6+(-6);
assign weight_bias7=in_buffer_weight7+(22);
assign weight_bias8=in_buffer_weight8+(-9);
assign weight_bias9=in_buffer_weight9+(59);
assign weight_bias10=in_buffer_weight10+(29);
assign weight_bias11=in_buffer_weight11+(-11);
assign weight_bias12=in_buffer_weight12+(-15);
assign weight_bias13=in_buffer_weight13+(-37);
assign weight_bias14=in_buffer_weight14+(52);
assign weight_bias15=in_buffer_weight15+(38);
assign weight_bias16=in_buffer_weight16+(37);
assign weight_bias17=in_buffer_weight17+(78);
assign weight_bias18=in_buffer_weight18+(-48);
assign weight_bias19=in_buffer_weight19+(-29);
assign weight_bias20=in_buffer_weight20+(8);
assign weight_bias21=in_buffer_weight21+(-21);
assign weight_bias22=in_buffer_weight22+(12);
assign weight_bias23=in_buffer_weight23+(77);
assign weight_bias24=in_buffer_weight24+(-10);
assign weight_bias25=in_buffer_weight25+(34);
assign weight_bias26=in_buffer_weight26+(17);
assign weight_bias27=in_buffer_weight27+(2);
assign weight_bias28=in_buffer_weight28+(55);
assign weight_bias29=in_buffer_weight29+(8);
assign weight_bias30=in_buffer_weight30+(-36);
assign weight_bias31=in_buffer_weight31+(23);
assign weight_bias32=in_buffer_weight32+(-29);
assign weight_bias33=in_buffer_weight33+(8);
assign weight_bias34=in_buffer_weight34+(0);
assign weight_bias35=in_buffer_weight35+(-25);
assign weight_bias36=in_buffer_weight36+(-27);
assign weight_bias37=in_buffer_weight37+(35);
assign weight_bias38=in_buffer_weight38+(-18);
assign weight_bias39=in_buffer_weight39+(50);
assign weight_bias40=in_buffer_weight40+(-28);
assign weight_bias41=in_buffer_weight41+(-2);
assign weight_bias42=in_buffer_weight42+(-47);
assign weight_bias43=in_buffer_weight43+(75);
assign weight_bias44=in_buffer_weight44+(51);
assign weight_bias45=in_buffer_weight45+(21);
assign weight_bias46=in_buffer_weight46+(-51);
assign weight_bias47=in_buffer_weight47+(14);
assign weight_bias48=in_buffer_weight48+(43);
assign weight_bias49=in_buffer_weight49+(-4);
assign weight_bias50=in_buffer_weight50+(55);
assign weight_bias51=in_buffer_weight51+(8);
assign weight_bias52=in_buffer_weight52+(19);
assign weight_bias53=in_buffer_weight53+(13);
assign weight_bias54=in_buffer_weight54+(94);
assign weight_bias55=in_buffer_weight55+(-9);
assign weight_bias56=in_buffer_weight56+(-13);
assign weight_bias57=in_buffer_weight57+(-21);
assign weight_bias58=in_buffer_weight58+(20);
assign weight_bias59=in_buffer_weight59+(5);
assign weight_bias60=in_buffer_weight60+(70);
assign weight_bias61=in_buffer_weight61+(-13);
assign weight_bias62=in_buffer_weight62+(28);
assign weight_bias63=in_buffer_weight63+(13);
wire signed [DATA_WIDTH-1:0]   bias_relu0;
wire signed [DATA_WIDTH-1:0]   bias_relu1;
wire signed [DATA_WIDTH-1:0]   bias_relu2;
wire signed [DATA_WIDTH-1:0]   bias_relu3;
wire signed [DATA_WIDTH-1:0]   bias_relu4;
wire signed [DATA_WIDTH-1:0]   bias_relu5;
wire signed [DATA_WIDTH-1:0]   bias_relu6;
wire signed [DATA_WIDTH-1:0]   bias_relu7;
wire signed [DATA_WIDTH-1:0]   bias_relu8;
wire signed [DATA_WIDTH-1:0]   bias_relu9;
wire signed [DATA_WIDTH-1:0]   bias_relu10;
wire signed [DATA_WIDTH-1:0]   bias_relu11;
wire signed [DATA_WIDTH-1:0]   bias_relu12;
wire signed [DATA_WIDTH-1:0]   bias_relu13;
wire signed [DATA_WIDTH-1:0]   bias_relu14;
wire signed [DATA_WIDTH-1:0]   bias_relu15;
wire signed [DATA_WIDTH-1:0]   bias_relu16;
wire signed [DATA_WIDTH-1:0]   bias_relu17;
wire signed [DATA_WIDTH-1:0]   bias_relu18;
wire signed [DATA_WIDTH-1:0]   bias_relu19;
wire signed [DATA_WIDTH-1:0]   bias_relu20;
wire signed [DATA_WIDTH-1:0]   bias_relu21;
wire signed [DATA_WIDTH-1:0]   bias_relu22;
wire signed [DATA_WIDTH-1:0]   bias_relu23;
wire signed [DATA_WIDTH-1:0]   bias_relu24;
wire signed [DATA_WIDTH-1:0]   bias_relu25;
wire signed [DATA_WIDTH-1:0]   bias_relu26;
wire signed [DATA_WIDTH-1:0]   bias_relu27;
wire signed [DATA_WIDTH-1:0]   bias_relu28;
wire signed [DATA_WIDTH-1:0]   bias_relu29;
wire signed [DATA_WIDTH-1:0]   bias_relu30;
wire signed [DATA_WIDTH-1:0]   bias_relu31;
wire signed [DATA_WIDTH-1:0]   bias_relu32;
wire signed [DATA_WIDTH-1:0]   bias_relu33;
wire signed [DATA_WIDTH-1:0]   bias_relu34;
wire signed [DATA_WIDTH-1:0]   bias_relu35;
wire signed [DATA_WIDTH-1:0]   bias_relu36;
wire signed [DATA_WIDTH-1:0]   bias_relu37;
wire signed [DATA_WIDTH-1:0]   bias_relu38;
wire signed [DATA_WIDTH-1:0]   bias_relu39;
wire signed [DATA_WIDTH-1:0]   bias_relu40;
wire signed [DATA_WIDTH-1:0]   bias_relu41;
wire signed [DATA_WIDTH-1:0]   bias_relu42;
wire signed [DATA_WIDTH-1:0]   bias_relu43;
wire signed [DATA_WIDTH-1:0]   bias_relu44;
wire signed [DATA_WIDTH-1:0]   bias_relu45;
wire signed [DATA_WIDTH-1:0]   bias_relu46;
wire signed [DATA_WIDTH-1:0]   bias_relu47;
wire signed [DATA_WIDTH-1:0]   bias_relu48;
wire signed [DATA_WIDTH-1:0]   bias_relu49;
wire signed [DATA_WIDTH-1:0]   bias_relu50;
wire signed [DATA_WIDTH-1:0]   bias_relu51;
wire signed [DATA_WIDTH-1:0]   bias_relu52;
wire signed [DATA_WIDTH-1:0]   bias_relu53;
wire signed [DATA_WIDTH-1:0]   bias_relu54;
wire signed [DATA_WIDTH-1:0]   bias_relu55;
wire signed [DATA_WIDTH-1:0]   bias_relu56;
wire signed [DATA_WIDTH-1:0]   bias_relu57;
wire signed [DATA_WIDTH-1:0]   bias_relu58;
wire signed [DATA_WIDTH-1:0]   bias_relu59;
wire signed [DATA_WIDTH-1:0]   bias_relu60;
wire signed [DATA_WIDTH-1:0]   bias_relu61;
wire signed [DATA_WIDTH-1:0]   bias_relu62;
wire signed [DATA_WIDTH-1:0]   bias_relu63;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign bias_relu32=(weight_bias32[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias32;
assign bias_relu33=(weight_bias33[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias33;
assign bias_relu34=(weight_bias34[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias34;
assign bias_relu35=(weight_bias35[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias35;
assign bias_relu36=(weight_bias36[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias36;
assign bias_relu37=(weight_bias37[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias37;
assign bias_relu38=(weight_bias38[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias38;
assign bias_relu39=(weight_bias39[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias39;
assign bias_relu40=(weight_bias40[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias40;
assign bias_relu41=(weight_bias41[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias41;
assign bias_relu42=(weight_bias42[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias42;
assign bias_relu43=(weight_bias43[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias43;
assign bias_relu44=(weight_bias44[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias44;
assign bias_relu45=(weight_bias45[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias45;
assign bias_relu46=(weight_bias46[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias46;
assign bias_relu47=(weight_bias47[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias47;
assign bias_relu48=(weight_bias48[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias48;
assign bias_relu49=(weight_bias49[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias49;
assign bias_relu50=(weight_bias50[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias50;
assign bias_relu51=(weight_bias51[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias51;
assign bias_relu52=(weight_bias52[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias52;
assign bias_relu53=(weight_bias53[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias53;
assign bias_relu54=(weight_bias54[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias54;
assign bias_relu55=(weight_bias55[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias55;
assign bias_relu56=(weight_bias56[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias56;
assign bias_relu57=(weight_bias57[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias57;
assign bias_relu58=(weight_bias58[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias58;
assign bias_relu59=(weight_bias59[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias59;
assign bias_relu60=(weight_bias60[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias60;
assign bias_relu61=(weight_bias61[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias61;
assign bias_relu62=(weight_bias62[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias62;
assign bias_relu63=(weight_bias63[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias63;
assign layer_out={bias_relu63,bias_relu62,bias_relu61,bias_relu60,bias_relu59,bias_relu58,bias_relu57,bias_relu56,bias_relu55,bias_relu54,bias_relu53,bias_relu52,bias_relu51,bias_relu50,bias_relu49,bias_relu48,bias_relu47,bias_relu46,bias_relu45,bias_relu44,bias_relu43,bias_relu42,bias_relu41,bias_relu40,bias_relu39,bias_relu38,bias_relu37,bias_relu36,bias_relu35,bias_relu34,bias_relu33,bias_relu32,bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule