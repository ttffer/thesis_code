module layer2_tcb_121x64x10
(
    input clk,
    input rst,
   input valid,
   output  reg ready,
    input [18*64-1:0]  layer_in,
    output [29*10-1:0]   layer_out
);
parameter DATA_WIDTH   =   29;
reg [DATA_WIDTH-1:0]    layer_in_buffer    [0:64-1];
integer i;
always@(posedge clk )
    begin
        if(rst)
            begin
                for(i=0;i<64;i=i+1)
                    begin
                        layer_in_buffer[i]<=0;
                    end
            end
        else
        begin
       layer_in_buffer[0]<=layer_in[17:0];
       layer_in_buffer[1]<=layer_in[35:18];
       layer_in_buffer[2]<=layer_in[53:36];
       layer_in_buffer[3]<=layer_in[71:54];
       layer_in_buffer[4]<=layer_in[89:72];
       layer_in_buffer[5]<=layer_in[107:90];
       layer_in_buffer[6]<=layer_in[125:108];
       layer_in_buffer[7]<=layer_in[143:126];
       layer_in_buffer[8]<=layer_in[161:144];
       layer_in_buffer[9]<=layer_in[179:162];
       layer_in_buffer[10]<=layer_in[197:180];
       layer_in_buffer[11]<=layer_in[215:198];
       layer_in_buffer[12]<=layer_in[233:216];
       layer_in_buffer[13]<=layer_in[251:234];
       layer_in_buffer[14]<=layer_in[269:252];
       layer_in_buffer[15]<=layer_in[287:270];
       layer_in_buffer[16]<=layer_in[305:288];
       layer_in_buffer[17]<=layer_in[323:306];
       layer_in_buffer[18]<=layer_in[341:324];
       layer_in_buffer[19]<=layer_in[359:342];
       layer_in_buffer[20]<=layer_in[377:360];
       layer_in_buffer[21]<=layer_in[395:378];
       layer_in_buffer[22]<=layer_in[413:396];
       layer_in_buffer[23]<=layer_in[431:414];
       layer_in_buffer[24]<=layer_in[449:432];
       layer_in_buffer[25]<=layer_in[467:450];
       layer_in_buffer[26]<=layer_in[485:468];
       layer_in_buffer[27]<=layer_in[503:486];
       layer_in_buffer[28]<=layer_in[521:504];
       layer_in_buffer[29]<=layer_in[539:522];
       layer_in_buffer[30]<=layer_in[557:540];
       layer_in_buffer[31]<=layer_in[575:558];
       layer_in_buffer[32]<=layer_in[593:576];
       layer_in_buffer[33]<=layer_in[611:594];
       layer_in_buffer[34]<=layer_in[629:612];
       layer_in_buffer[35]<=layer_in[647:630];
       layer_in_buffer[36]<=layer_in[665:648];
       layer_in_buffer[37]<=layer_in[683:666];
       layer_in_buffer[38]<=layer_in[701:684];
       layer_in_buffer[39]<=layer_in[719:702];
       layer_in_buffer[40]<=layer_in[737:720];
       layer_in_buffer[41]<=layer_in[755:738];
       layer_in_buffer[42]<=layer_in[773:756];
       layer_in_buffer[43]<=layer_in[791:774];
       layer_in_buffer[44]<=layer_in[809:792];
       layer_in_buffer[45]<=layer_in[827:810];
       layer_in_buffer[46]<=layer_in[845:828];
       layer_in_buffer[47]<=layer_in[863:846];
       layer_in_buffer[48]<=layer_in[881:864];
       layer_in_buffer[49]<=layer_in[899:882];
       layer_in_buffer[50]<=layer_in[917:900];
       layer_in_buffer[51]<=layer_in[935:918];
       layer_in_buffer[52]<=layer_in[953:936];
       layer_in_buffer[53]<=layer_in[971:954];
       layer_in_buffer[54]<=layer_in[989:972];
       layer_in_buffer[55]<=layer_in[1007:990];
       layer_in_buffer[56]<=layer_in[1025:1008];
       layer_in_buffer[57]<=layer_in[1043:1026];
       layer_in_buffer[58]<=layer_in[1061:1044];
       layer_in_buffer[59]<=layer_in[1079:1062];
       layer_in_buffer[60]<=layer_in[1097:1080];
       layer_in_buffer[61]<=layer_in[1115:1098];
       layer_in_buffer[62]<=layer_in[1133:1116];
       layer_in_buffer[63]<=layer_in[1151:1134];
        end
   end

wire [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0-(0-(layer_in_buffer[0]<<1)-(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<7))+(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<6))-(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<6))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<6))+(0-(layer_in_buffer[6]<<0)-(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<6))+(0-(layer_in_buffer[7]<<0)-(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<6))-(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6))+(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6))-(0-(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<6))-(0-(layer_in_buffer[13]<<1)-(layer_in_buffer[13]<<3)+(layer_in_buffer[13]<<7))+(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<6))+(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<6))+(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<6))+(0-(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<6))-(0-(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<6))+(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<6))-(0-(layer_in_buffer[24]<<0)-(layer_in_buffer[24]<<2)+(layer_in_buffer[24]<<6))-(0-(layer_in_buffer[25]<<0)-(layer_in_buffer[25]<<2)+(layer_in_buffer[25]<<6))+(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))-(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<6))+(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<6))+(0-(layer_in_buffer[34]<<0)-(layer_in_buffer[34]<<2)+(layer_in_buffer[34]<<6))+(0-(layer_in_buffer[38]<<0)-(layer_in_buffer[38]<<2)+(layer_in_buffer[38]<<6))-(0-(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<2)+(layer_in_buffer[40]<<6))+(0-(layer_in_buffer[41]<<0)-(layer_in_buffer[41]<<2)+(layer_in_buffer[41]<<6))-(0-(layer_in_buffer[43]<<0)-(layer_in_buffer[43]<<2)+(layer_in_buffer[43]<<6))-(0-(layer_in_buffer[44]<<1)-(layer_in_buffer[44]<<3)+(layer_in_buffer[44]<<7))+(0-(layer_in_buffer[45]<<0)-(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6))+(0-(layer_in_buffer[46]<<0)-(layer_in_buffer[46]<<2)+(layer_in_buffer[46]<<6))+(0-(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<6))-(0-(layer_in_buffer[48]<<1)-(layer_in_buffer[48]<<3)+(layer_in_buffer[48]<<7))-(0-(layer_in_buffer[52]<<0)-(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<6))-(0+(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<4)+(layer_in_buffer[54]<<6)+(layer_in_buffer[54]<<7))-(0-(layer_in_buffer[55]<<0)-(layer_in_buffer[55]<<2)+(layer_in_buffer[55]<<6))+(0-(layer_in_buffer[56]<<1)-(layer_in_buffer[56]<<3)+(layer_in_buffer[56]<<7))+(0-(layer_in_buffer[58]<<0)-(layer_in_buffer[58]<<2)+(layer_in_buffer[58]<<6))+(0-(layer_in_buffer[59]<<0)-(layer_in_buffer[59]<<2)+(layer_in_buffer[59]<<6))-(0+(layer_in_buffer[61]<<0)-(layer_in_buffer[61]<<4)+(layer_in_buffer[61]<<6)+(layer_in_buffer[61]<<7))-(0-(layer_in_buffer[62]<<1)-(layer_in_buffer[62]<<3)+(layer_in_buffer[62]<<7));
wire [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0+(0-(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<6))+(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<6))+(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<6))-(0-(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6))-(0-(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<6))+(0-(layer_in_buffer[6]<<0)-(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<6))-(0-(layer_in_buffer[7]<<0)-(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<6))-(0-(layer_in_buffer[8]<<1)-(layer_in_buffer[8]<<3)+(layer_in_buffer[8]<<7))+(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6))-(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<6))-(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6))+(0+(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<6)+(layer_in_buffer[14]<<7))-(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<6))-(0-(layer_in_buffer[16]<<1)-(layer_in_buffer[16]<<3)+(layer_in_buffer[16]<<7))+(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<6))+(0-(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6))-(0-(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<6))+(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<6))-(0-(layer_in_buffer[24]<<1)-(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<7))-(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))-(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))-(0-(layer_in_buffer[29]<<0)-(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<6))-(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<6))-(0-(layer_in_buffer[34]<<1)-(layer_in_buffer[34]<<3)+(layer_in_buffer[34]<<7))+(0-(layer_in_buffer[35]<<0)-(layer_in_buffer[35]<<2)+(layer_in_buffer[35]<<6))+(0-(layer_in_buffer[36]<<0)-(layer_in_buffer[36]<<2)+(layer_in_buffer[36]<<6))-(0-(layer_in_buffer[37]<<1)-(layer_in_buffer[37]<<3)+(layer_in_buffer[37]<<7))-(0-(layer_in_buffer[38]<<1)-(layer_in_buffer[38]<<3)+(layer_in_buffer[38]<<7))-(0-(layer_in_buffer[40]<<1)-(layer_in_buffer[40]<<3)+(layer_in_buffer[40]<<7))-(0-(layer_in_buffer[41]<<0)-(layer_in_buffer[41]<<2)+(layer_in_buffer[41]<<6))+(0-(layer_in_buffer[42]<<0)-(layer_in_buffer[42]<<2)+(layer_in_buffer[42]<<6))-(0-(layer_in_buffer[45]<<1)-(layer_in_buffer[45]<<3)+(layer_in_buffer[45]<<7))-(0-(layer_in_buffer[46]<<0)-(layer_in_buffer[46]<<2)+(layer_in_buffer[46]<<6))+(0-(layer_in_buffer[48]<<1)-(layer_in_buffer[48]<<3)+(layer_in_buffer[48]<<7))-(0-(layer_in_buffer[50]<<0)-(layer_in_buffer[50]<<2)+(layer_in_buffer[50]<<6))+(0-(layer_in_buffer[51]<<0)-(layer_in_buffer[51]<<2)+(layer_in_buffer[51]<<6))+(0-(layer_in_buffer[52]<<0)-(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<6))-(0-(layer_in_buffer[53]<<1)-(layer_in_buffer[53]<<3)+(layer_in_buffer[53]<<7))+(0-(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<6))+(0-(layer_in_buffer[56]<<0)-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<6))+(0+(layer_in_buffer[58]<<0)-(layer_in_buffer[58]<<4)+(layer_in_buffer[58]<<6)+(layer_in_buffer[58]<<7))-(0-(layer_in_buffer[60]<<0)-(layer_in_buffer[60]<<2)+(layer_in_buffer[60]<<6))-(0-(layer_in_buffer[61]<<1)-(layer_in_buffer[61]<<3)+(layer_in_buffer[61]<<7))+(0-(layer_in_buffer[62]<<0)-(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0+(0-(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<6))+(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<6))+(0-(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<6))+(0-(layer_in_buffer[5]<<1)-(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<7))-(0-(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<6))+(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<6))+(0-(layer_in_buffer[13]<<0)-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<6))-(0-(layer_in_buffer[14]<<2)-(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<8))-(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<6))-(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<6))+(0-(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<6))-(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<6))+(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<6))+(0-(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6))+(0-(layer_in_buffer[25]<<1)-(layer_in_buffer[25]<<3)+(layer_in_buffer[25]<<7))-(0-(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<2)+(layer_in_buffer[26]<<6))+(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))+(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))+(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<6))-(0-(layer_in_buffer[34]<<0)-(layer_in_buffer[34]<<2)+(layer_in_buffer[34]<<6))-(0-(layer_in_buffer[35]<<1)-(layer_in_buffer[35]<<3)+(layer_in_buffer[35]<<7))+(0-(layer_in_buffer[39]<<0)-(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<6))-(0-(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<2)+(layer_in_buffer[40]<<6))-(0-(layer_in_buffer[42]<<2)-(layer_in_buffer[42]<<4)+(layer_in_buffer[42]<<8))-(0-(layer_in_buffer[43]<<0)-(layer_in_buffer[43]<<2)+(layer_in_buffer[43]<<6))-(0-(layer_in_buffer[45]<<0)-(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6))+(0-(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<6))-(0-(layer_in_buffer[48]<<0)-(layer_in_buffer[48]<<2)+(layer_in_buffer[48]<<6))+(0-(layer_in_buffer[49]<<0)-(layer_in_buffer[49]<<2)+(layer_in_buffer[49]<<6))+(0-(layer_in_buffer[51]<<0)-(layer_in_buffer[51]<<2)+(layer_in_buffer[51]<<6))+(0-(layer_in_buffer[53]<<0)-(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<6))-(0-(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<6))+(0-(layer_in_buffer[56]<<0)-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<6))+(0-(layer_in_buffer[58]<<0)-(layer_in_buffer[58]<<2)+(layer_in_buffer[58]<<6))-(0-(layer_in_buffer[61]<<0)-(layer_in_buffer[61]<<2)+(layer_in_buffer[61]<<6))+(0-(layer_in_buffer[63]<<0)-(layer_in_buffer[63]<<2)+(layer_in_buffer[63]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0-(0-(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<7))-(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<6))+(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<6))+(0-(layer_in_buffer[6]<<0)-(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<6))-(0-(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<6))-(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6))-(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<6))+(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6))-(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<6))+(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<6))-(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<6))+(0-(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<6))+(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<6))+(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<6))+(0-(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6))-(0-(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<6))-(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<6))+(0-(layer_in_buffer[24]<<0)-(layer_in_buffer[24]<<2)+(layer_in_buffer[24]<<6))-(0-(layer_in_buffer[25]<<0)-(layer_in_buffer[25]<<2)+(layer_in_buffer[25]<<6))-(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))+(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))-(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<6))-(0+(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<6)+(layer_in_buffer[31]<<7))+(0-(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<2)+(layer_in_buffer[33]<<6))+(0-(layer_in_buffer[35]<<0)-(layer_in_buffer[35]<<2)+(layer_in_buffer[35]<<6))-(0+(layer_in_buffer[36]<<0)-(layer_in_buffer[36]<<4)+(layer_in_buffer[36]<<6)+(layer_in_buffer[36]<<7))-(0-(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<2)+(layer_in_buffer[37]<<6))+(0-(layer_in_buffer[39]<<0)-(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<6))-(0-(layer_in_buffer[42]<<1)-(layer_in_buffer[42]<<3)+(layer_in_buffer[42]<<7))+(0-(layer_in_buffer[43]<<0)-(layer_in_buffer[43]<<2)+(layer_in_buffer[43]<<6))+(0-(layer_in_buffer[44]<<0)-(layer_in_buffer[44]<<2)+(layer_in_buffer[44]<<6))-(0-(layer_in_buffer[45]<<1)-(layer_in_buffer[45]<<3)+(layer_in_buffer[45]<<7))+(0-(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<6))+(0-(layer_in_buffer[51]<<0)-(layer_in_buffer[51]<<2)+(layer_in_buffer[51]<<6))-(0-(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<6))-(0-(layer_in_buffer[56]<<0)-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<6))-(0-(layer_in_buffer[58]<<1)-(layer_in_buffer[58]<<3)+(layer_in_buffer[58]<<7))+(0-(layer_in_buffer[59]<<0)-(layer_in_buffer[59]<<2)+(layer_in_buffer[59]<<6))+(0-(layer_in_buffer[60]<<0)-(layer_in_buffer[60]<<2)+(layer_in_buffer[60]<<6))+(0-(layer_in_buffer[61]<<1)-(layer_in_buffer[61]<<3)+(layer_in_buffer[61]<<7))-(0-(layer_in_buffer[63]<<0)-(layer_in_buffer[63]<<2)+(layer_in_buffer[63]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0+(0-(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<6))+(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<6))-(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<6))+(0-(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<6))-(0-(layer_in_buffer[6]<<2)-(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<8))+(0-(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<6))-(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6))+(0-(layer_in_buffer[13]<<0)-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<6))+(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<6))-(0+(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<4)+(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<7))-(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<6))-(0-(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<4)+(layer_in_buffer[19]<<8))-(0-(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6))-(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<6))-(0-(layer_in_buffer[25]<<0)-(layer_in_buffer[25]<<2)+(layer_in_buffer[25]<<6))-(0-(layer_in_buffer[27]<<1)-(layer_in_buffer[27]<<3)+(layer_in_buffer[27]<<7))-(0+(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<4)+(layer_in_buffer[28]<<6)+(layer_in_buffer[28]<<7))+(0-(layer_in_buffer[29]<<0)-(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<6))+(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<6))+(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<6))-(0-(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<2)+(layer_in_buffer[33]<<6))+(0-(layer_in_buffer[35]<<0)-(layer_in_buffer[35]<<2)+(layer_in_buffer[35]<<6))-(0-(layer_in_buffer[36]<<0)-(layer_in_buffer[36]<<2)+(layer_in_buffer[36]<<6))+(0-(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<2)+(layer_in_buffer[37]<<6))+(0-(layer_in_buffer[39]<<0)-(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<6))+(0-(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<2)+(layer_in_buffer[40]<<6))-(0-(layer_in_buffer[41]<<0)-(layer_in_buffer[41]<<2)+(layer_in_buffer[41]<<6))-(0-(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<6))-(0-(layer_in_buffer[48]<<0)-(layer_in_buffer[48]<<2)+(layer_in_buffer[48]<<6))-(0+(layer_in_buffer[49]<<0)-(layer_in_buffer[49]<<4)+(layer_in_buffer[49]<<6)+(layer_in_buffer[49]<<7))-(0-(layer_in_buffer[52]<<0)-(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<6))+(0-(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<6))-(0-(layer_in_buffer[55]<<2)-(layer_in_buffer[55]<<4)+(layer_in_buffer[55]<<8))+(0-(layer_in_buffer[59]<<0)-(layer_in_buffer[59]<<2)+(layer_in_buffer[59]<<6))-(0-(layer_in_buffer[60]<<1)-(layer_in_buffer[60]<<3)+(layer_in_buffer[60]<<7))+(0-(layer_in_buffer[61]<<0)-(layer_in_buffer[61]<<2)+(layer_in_buffer[61]<<6))+(0-(layer_in_buffer[63]<<0)-(layer_in_buffer[63]<<2)+(layer_in_buffer[63]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0+(0-(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<6))-(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<6))+(0-(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<6))-(0-(layer_in_buffer[6]<<0)-(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<6))-(0-(layer_in_buffer[7]<<1)-(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<7))+(0-(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<6))+(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6))-(0+(layer_in_buffer[13]<<0)-(layer_in_buffer[13]<<4)+(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<7))+(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<6))-(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<6))-(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<6))-(0-(layer_in_buffer[17]<<1)-(layer_in_buffer[17]<<3)+(layer_in_buffer[17]<<7))+(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<6))-(0-(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6))+(0-(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<6))+(0-(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<2)+(layer_in_buffer[26]<<6))+(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))-(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))+(0-(layer_in_buffer[29]<<0)-(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<6))-(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<6))-(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<6))-(0-(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<2)+(layer_in_buffer[33]<<6))+(0-(layer_in_buffer[37]<<1)-(layer_in_buffer[37]<<3)+(layer_in_buffer[37]<<7))+(0-(layer_in_buffer[38]<<0)-(layer_in_buffer[38]<<2)+(layer_in_buffer[38]<<6))-(0-(layer_in_buffer[39]<<2)-(layer_in_buffer[39]<<4)+(layer_in_buffer[39]<<8))+(0-(layer_in_buffer[42]<<0)-(layer_in_buffer[42]<<2)+(layer_in_buffer[42]<<6))+(0-(layer_in_buffer[44]<<0)-(layer_in_buffer[44]<<2)+(layer_in_buffer[44]<<6))+(0-(layer_in_buffer[45]<<0)-(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6))+(0-(layer_in_buffer[49]<<0)-(layer_in_buffer[49]<<2)+(layer_in_buffer[49]<<6))-(0-(layer_in_buffer[51]<<2)-(layer_in_buffer[51]<<4)+(layer_in_buffer[51]<<8))+(0-(layer_in_buffer[52]<<0)-(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<6))-(0-(layer_in_buffer[53]<<0)-(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<6))+(0-(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<6))+(0-(layer_in_buffer[55]<<1)-(layer_in_buffer[55]<<3)+(layer_in_buffer[55]<<7))-(0-(layer_in_buffer[56]<<0)+(layer_in_buffer[56]<<3)+(layer_in_buffer[56]<<5)+(layer_in_buffer[56]<<8))+(0-(layer_in_buffer[58]<<0)-(layer_in_buffer[58]<<2)+(layer_in_buffer[58]<<6))+(0-(layer_in_buffer[61]<<0)-(layer_in_buffer[61]<<2)+(layer_in_buffer[61]<<6))+(0-(layer_in_buffer[62]<<0)-(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<6))-(0-(layer_in_buffer[63]<<0)-(layer_in_buffer[63]<<2)+(layer_in_buffer[63]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0+(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<6))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<6))+(0-(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<6))-(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6))+(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<6))+(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6))+(0-(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<6))+(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<6))+(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<6))-(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<6))-(0-(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6))+(0-(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<6))-(0-(layer_in_buffer[24]<<1)-(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<7))-(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))+(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))-(0+(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<4)+(layer_in_buffer[33]<<6)+(layer_in_buffer[33]<<7))-(0-(layer_in_buffer[34]<<0)-(layer_in_buffer[34]<<2)+(layer_in_buffer[34]<<6))+(0-(layer_in_buffer[36]<<0)-(layer_in_buffer[36]<<2)+(layer_in_buffer[36]<<6))-(0+(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<4)+(layer_in_buffer[37]<<6)+(layer_in_buffer[37]<<7))-(0-(layer_in_buffer[38]<<0)-(layer_in_buffer[38]<<2)+(layer_in_buffer[38]<<6))-(0-(layer_in_buffer[39]<<1)-(layer_in_buffer[39]<<3)+(layer_in_buffer[39]<<7))+(0-(layer_in_buffer[42]<<0)-(layer_in_buffer[42]<<2)+(layer_in_buffer[42]<<6))-(0-(layer_in_buffer[43]<<1)-(layer_in_buffer[43]<<3)+(layer_in_buffer[43]<<7))-(0+(layer_in_buffer[44]<<0)-(layer_in_buffer[44]<<4)+(layer_in_buffer[44]<<6)+(layer_in_buffer[44]<<7))+(0-(layer_in_buffer[45]<<0)-(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6))+(0-(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<6))-(0-(layer_in_buffer[49]<<0)-(layer_in_buffer[49]<<2)+(layer_in_buffer[49]<<6))-(0+(layer_in_buffer[51]<<0)-(layer_in_buffer[51]<<4)+(layer_in_buffer[51]<<6)+(layer_in_buffer[51]<<7))+(0-(layer_in_buffer[53]<<0)-(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<6))-(0-(layer_in_buffer[54]<<1)-(layer_in_buffer[54]<<3)+(layer_in_buffer[54]<<7))+(0-(layer_in_buffer[55]<<0)-(layer_in_buffer[55]<<2)+(layer_in_buffer[55]<<6))+(0-(layer_in_buffer[56]<<0)-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<6))+(0-(layer_in_buffer[60]<<0)-(layer_in_buffer[60]<<2)+(layer_in_buffer[60]<<6))-(0+(layer_in_buffer[61]<<0)-(layer_in_buffer[61]<<4)+(layer_in_buffer[61]<<6)+(layer_in_buffer[61]<<7))-(0-(layer_in_buffer[62]<<0)-(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<6))+(0-(layer_in_buffer[63]<<0)-(layer_in_buffer[63]<<2)+(layer_in_buffer[63]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0-(0-(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<6))-(0-(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<7))+(0+(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<4)+(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<7))-(0-(layer_in_buffer[3]<<1)-(layer_in_buffer[3]<<3)+(layer_in_buffer[3]<<7))+(0-(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<6))+(0-(layer_in_buffer[7]<<0)-(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<6))+(0-(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<6))+(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6))-(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<6))-(0-(layer_in_buffer[11]<<1)-(layer_in_buffer[11]<<3)+(layer_in_buffer[11]<<7))-(0-(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<6))+(0-(layer_in_buffer[13]<<0)-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<6))-(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<6))+(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<6))-(0-(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6))+(0-(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<6))-(0-(layer_in_buffer[22]<<1)-(layer_in_buffer[22]<<3)+(layer_in_buffer[22]<<7))+(0-(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<2)+(layer_in_buffer[26]<<6))+(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))+(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))-(0-(layer_in_buffer[29]<<0)-(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<6))-(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<6))+(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<6))+(0-(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<2)+(layer_in_buffer[33]<<6))+(0-(layer_in_buffer[34]<<0)-(layer_in_buffer[34]<<2)+(layer_in_buffer[34]<<6))+(0-(layer_in_buffer[35]<<1)-(layer_in_buffer[35]<<3)+(layer_in_buffer[35]<<7))+(0-(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<2)+(layer_in_buffer[37]<<6))+(0-(layer_in_buffer[39]<<0)-(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<6))+(0-(layer_in_buffer[41]<<0)-(layer_in_buffer[41]<<2)+(layer_in_buffer[41]<<6))-(0-(layer_in_buffer[45]<<0)-(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6))-(0-(layer_in_buffer[46]<<0)-(layer_in_buffer[46]<<2)+(layer_in_buffer[46]<<6))+(0-(layer_in_buffer[48]<<0)-(layer_in_buffer[48]<<2)+(layer_in_buffer[48]<<6))-(0-(layer_in_buffer[49]<<0)-(layer_in_buffer[49]<<2)+(layer_in_buffer[49]<<6))-(0-(layer_in_buffer[50]<<1)-(layer_in_buffer[50]<<3)+(layer_in_buffer[50]<<7))-(0-(layer_in_buffer[52]<<0)-(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<6))-(0-(layer_in_buffer[53]<<0)-(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<6))+(0-(layer_in_buffer[56]<<0)-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<6))-(0-(layer_in_buffer[58]<<1)-(layer_in_buffer[58]<<3)+(layer_in_buffer[58]<<7))-(0-(layer_in_buffer[59]<<0)-(layer_in_buffer[59]<<2)+(layer_in_buffer[59]<<6))-(0-(layer_in_buffer[60]<<1)-(layer_in_buffer[60]<<3)+(layer_in_buffer[60]<<7))+(0-(layer_in_buffer[61]<<0)-(layer_in_buffer[61]<<2)+(layer_in_buffer[61]<<6))-(0-(layer_in_buffer[63]<<0)-(layer_in_buffer[63]<<2)+(layer_in_buffer[63]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0-(0-(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<7))-(0-(layer_in_buffer[2]<<1)-(layer_in_buffer[2]<<3)+(layer_in_buffer[2]<<7))+(0-(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6))-(0+(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<6)+(layer_in_buffer[5]<<7))+(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<6))-(0-(layer_in_buffer[14]<<1)-(layer_in_buffer[14]<<3)+(layer_in_buffer[14]<<7))-(0-(layer_in_buffer[15]<<1)-(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<7))+(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<6))-(0-(layer_in_buffer[19]<<1)-(layer_in_buffer[19]<<3)+(layer_in_buffer[19]<<7))+(0-(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<6))+(0-(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<6))+(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<6))+(0-(layer_in_buffer[25]<<0)-(layer_in_buffer[25]<<2)+(layer_in_buffer[25]<<6))-(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6))-(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))-(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<6))-(0-(layer_in_buffer[35]<<1)-(layer_in_buffer[35]<<3)+(layer_in_buffer[35]<<7))+(0-(layer_in_buffer[36]<<0)-(layer_in_buffer[36]<<2)+(layer_in_buffer[36]<<6))-(0-(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<2)+(layer_in_buffer[37]<<6))+(0-(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<2)+(layer_in_buffer[40]<<6))+(0-(layer_in_buffer[46]<<0)-(layer_in_buffer[46]<<2)+(layer_in_buffer[46]<<6))-(0-(layer_in_buffer[47]<<1)-(layer_in_buffer[47]<<3)+(layer_in_buffer[47]<<7))-(0-(layer_in_buffer[48]<<1)-(layer_in_buffer[48]<<3)+(layer_in_buffer[48]<<7))+(0-(layer_in_buffer[50]<<0)-(layer_in_buffer[50]<<2)+(layer_in_buffer[50]<<6))+(0-(layer_in_buffer[52]<<0)-(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<6))-(0-(layer_in_buffer[53]<<0)-(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<6))-(0-(layer_in_buffer[56]<<0)-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<6))-(0-(layer_in_buffer[58]<<1)-(layer_in_buffer[58]<<3)+(layer_in_buffer[58]<<7))+(0-(layer_in_buffer[60]<<0)-(layer_in_buffer[60]<<2)+(layer_in_buffer[60]<<6))-(0-(layer_in_buffer[61]<<0)-(layer_in_buffer[61]<<2)+(layer_in_buffer[61]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0-(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<6)+(layer_in_buffer[0]<<7))+(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<6))-(0-(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<3)+(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<8))+(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<6))-(0+(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<6)+(layer_in_buffer[5]<<7))+(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6))-(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<6))-(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6))+(0-(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<6))-(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<6))-(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<6))+(0-(layer_in_buffer[24]<<0)-(layer_in_buffer[24]<<2)+(layer_in_buffer[24]<<6))-(0-(layer_in_buffer[25]<<2)-(layer_in_buffer[25]<<4)+(layer_in_buffer[25]<<8))-(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<6))+(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<6))+(0-(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<2)+(layer_in_buffer[33]<<6))-(0-(layer_in_buffer[36]<<2)-(layer_in_buffer[36]<<4)+(layer_in_buffer[36]<<8))+(0-(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<2)+(layer_in_buffer[37]<<6))+(0-(layer_in_buffer[42]<<0)-(layer_in_buffer[42]<<2)+(layer_in_buffer[42]<<6))-(0-(layer_in_buffer[43]<<0)-(layer_in_buffer[43]<<2)+(layer_in_buffer[43]<<6))+(0-(layer_in_buffer[45]<<0)-(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6))-(0+(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<4)+(layer_in_buffer[47]<<6)+(layer_in_buffer[47]<<7))-(0-(layer_in_buffer[49]<<1)-(layer_in_buffer[49]<<3)+(layer_in_buffer[49]<<7))+(0-(layer_in_buffer[51]<<0)-(layer_in_buffer[51]<<2)+(layer_in_buffer[51]<<6))+(0-(layer_in_buffer[53]<<0)-(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<6))+(0-(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<6))-(0-(layer_in_buffer[55]<<0)-(layer_in_buffer[55]<<2)+(layer_in_buffer[55]<<6))+(0-(layer_in_buffer[56]<<0)-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<6))-(0+(layer_in_buffer[58]<<0)-(layer_in_buffer[58]<<4)+(layer_in_buffer[58]<<6)+(layer_in_buffer[58]<<7))-(0-(layer_in_buffer[59]<<1)-(layer_in_buffer[59]<<3)+(layer_in_buffer[59]<<7))+(0-(layer_in_buffer[60]<<0)-(layer_in_buffer[60]<<2)+(layer_in_buffer[60]<<6))-(0-(layer_in_buffer[62]<<0)-(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<6));
wire [DATA_WIDTH-1:0]   weight_bias0;
assign weight_bias0=in_buffer_weight0+(0);
wire [DATA_WIDTH-1:0]   weight_bias1;
assign weight_bias1=in_buffer_weight1+(0);
wire [DATA_WIDTH-1:0]   weight_bias2;
assign weight_bias2=in_buffer_weight2+(0);
wire [DATA_WIDTH-1:0]   weight_bias3;
assign weight_bias3=in_buffer_weight3+(0);
wire [DATA_WIDTH-1:0]   weight_bias4;
assign weight_bias4=in_buffer_weight4+(0);
wire [DATA_WIDTH-1:0]   weight_bias5;
assign weight_bias5=in_buffer_weight5+(59);
wire [DATA_WIDTH-1:0]   weight_bias6;
assign weight_bias6=in_buffer_weight6+(0);
wire [DATA_WIDTH-1:0]   weight_bias7;
assign weight_bias7=in_buffer_weight7+(0);
wire [DATA_WIDTH-1:0]   weight_bias8;
assign weight_bias8=in_buffer_weight8+(0);
wire [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias9=in_buffer_weight9+(0);
assign layer_out={
            weight_bias9,
            weight_bias8,
            weight_bias7,
            weight_bias6,
            weight_bias5,
            weight_bias4,
            weight_bias3,
            weight_bias2,
            weight_bias1,
            weight_bias0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule
