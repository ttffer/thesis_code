module barrett_n13(input [5:0] codeword,output [2:0]q,output [3:0]r,output error,output[5:0] receive);
    wire[9:0]q_temp;
    wire[4:0]r_temp;
    assign q_temp=codeword*4'd9>>7;
    assign r_temp=codeword-q_temp*4'd13;
    assign q=r_temp<4'd13 ? q_temp:q_temp+1'b1;
    assign r=r_temp<4'd13 ? r_temp:r_temp-4'd13;
    assign error = r|4'b0 ? 1'b1:1'b0;
    assign receive = codeword;
endmodule