`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/23/2022 04:22:55 AM
// Design Name: 
// Module Name: n13sys6x6_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module n13sys6x6_testbench(

    );
    
    reg [5:0]word0,word1,word2,word3,word4,word5,word6,word7,word8,word9,word10,word11,word12,word13,word14,word15,word16,word17,word18,word19,word20,word21,word22,word23,word24,word25,word26,word27,word28,word29,word30,word31,word32,word33,word34,word35;
    wire [2:0]d_word0,d_word1,d_word2,d_word3,d_word4,d_word5,d_word6,d_word7,d_word8,d_word9,d_word10,d_word11,d_word12,d_word13,d_word14,d_word15,d_word16,d_word17,d_word18,d_word19,d_word20,d_word21,d_word22,d_word23,d_word24,d_word25,d_word26,d_word27,d_word28,d_word29,d_word30,d_word31,d_word32,d_word33,d_word34,d_word35;
    n13sys_6x6 DUT_n13(.IN0(word0),.IN1(word1),.IN2(word2),.IN3(word3),.IN4(word4),.IN5(word5),.IN6(word6),.IN7(word7),.IN8(word8),.IN9(word9),.IN10(word10),.IN11(word11),.IN12(word12),.IN13(word13),.IN14(word14),.IN15(word15),.IN16(word16),.IN17(word17),.IN18(word18),.IN19(word19),.IN20(word20),.IN21(word21),.IN22(word22),.IN23(word23),.IN24(word24),.IN25(word25),.IN26(word26),.IN27(word27),.IN28(word28),.IN29(word29),.IN30(word30),.IN31(word31),.IN32(word32),.IN33(word33),.IN34(word34),.IN35(word35)
                    ,.OUT0(d_word0),.OUT1(d_word1),.OUT2(d_word2),.OUT3(d_word3),.OUT4(d_word4),.OUT5(d_word5),.OUT6(d_word6),.OUT7(d_word7),.OUT8(d_word8),.OUT9(d_word9),.OUT10(d_word10),.OUT11(d_word11),.OUT12(d_word12),.OUT13(d_word13),.OUT14(d_word14),.OUT15(d_word15),.OUT16(d_word16),.OUT17(d_word17),.OUT18(d_word18),.OUT19(d_word19),.OUT20(d_word20),.OUT21(d_word21),.OUT22(d_word22),.OUT23(d_word23),.OUT24(d_word24),.OUT25(d_word25),.OUT26(d_word26),.OUT27(d_word27),.OUT28(d_word28),.OUT29(d_word29),.OUT30(d_word30),.OUT31(d_word31),.OUT32(d_word32),.OUT33(d_word33),.OUT34(d_word34),.OUT35(d_word35));
    
    initial begin 
    word0='d0;word1='d0;word2='d0;word3='d0;word4='d0;word5='d0;word6='d0;word7='d0;word8='d0;word9='d0;word10='d0;word11='d0;word12='d0;word13='d0;word14='d0;word15='d0;word16='d0;word17='d0;word18='d0;word19='d0;word20='d0;word21='d0;word22='d0;word23='d0;word24='d0;word25='d0;word26='d0;word27='d0;word28='d0;word29='d0;word30='d0;word31='d0;word32='d0;word33='d0;word34='d0;word35='d0;
    #10 word0='d13;
#10 word0='d26;
#10 word0='d39;
#10 word0='d52;
#10 word0='d1;
#10 word0='d0;#10 word1='d1;
#10 word1='d0;#10 word2='d1;
#10 word2='d0;#10 word3='d1;
#10 word3='d0;#10 word4='d1;
#10 word4='d0;#10 word5='d1;
#10 word5='d0;#10 word6='d1;
#10 word6='d0;#10 word7='d1;
#10 word7='d0;#10 word8='d1;
#10 word8='d0;#10 word9='d1;
#10 word9='d0;#10 word10='d1;
#10 word10='d0;#10 word11='d1;
#10 word11='d0;#10 word12='d1;
#10 word12='d0;#10 word13='d1;
#10 word13='d0;#10 word14='d1;
#10 word14='d0;#10 word15='d1;
#10 word15='d0;#10 word16='d1;
#10 word16='d0;#10 word17='d1;
#10 word17='d0;#10 word18='d1;
#10 word18='d0;#10 word19='d1;
#10 word19='d0;#10 word20='d1;
#10 word20='d0;#10 word21='d1;
#10 word21='d0;#10 word22='d1;
#10 word22='d0;#10 word23='d1;
#10 word23='d0;#10 word24='d1;
#10 word24='d0;#10 word25='d1;
#10 word25='d0;#10 word26='d1;
#10 word26='d0;#10 word27='d1;
#10 word27='d0;#10 word28='d1;
#10 word28='d0;#10 word29='d1;
#10 word29='d0;#10 word30='d1;
#10 word30='d0;#10 word31='d1;
#10 word31='d0;#10 word32='d1;
#10 word32='d0;#10 word33='d1;
#10 word33='d0;#10 word34='d1;
#10 word34='d0;#10 word35='d1;
#10 word35='d0;#10 word0='d2;
#10 word0='d0;#10 word1='d2;
#10 word1='d0;#10 word2='d2;
#10 word2='d0;#10 word3='d2;
#10 word3='d0;#10 word4='d2;
#10 word4='d0;#10 word5='d2;
#10 word5='d0;#10 word6='d2;
#10 word6='d0;#10 word7='d2;
#10 word7='d0;#10 word8='d2;
#10 word8='d0;#10 word9='d2;
#10 word9='d0;#10 word10='d2;
#10 word10='d0;#10 word11='d2;
#10 word11='d0;#10 word12='d2;
#10 word12='d0;#10 word13='d2;
#10 word13='d0;#10 word14='d2;
#10 word14='d0;#10 word15='d2;
#10 word15='d0;#10 word16='d2;
#10 word16='d0;#10 word17='d2;
#10 word17='d0;#10 word18='d2;
#10 word18='d0;#10 word19='d2;
#10 word19='d0;#10 word20='d2;
#10 word20='d0;#10 word21='d2;
#10 word21='d0;#10 word22='d2;
#10 word22='d0;#10 word23='d2;
#10 word23='d0;#10 word24='d2;
#10 word24='d0;#10 word25='d2;
#10 word25='d0;#10 word26='d2;
#10 word26='d0;#10 word27='d2;
#10 word27='d0;#10 word28='d2;
#10 word28='d0;#10 word29='d2;
#10 word29='d0;#10 word30='d2;
#10 word30='d0;#10 word31='d2;
#10 word31='d0;#10 word32='d2;
#10 word32='d0;#10 word33='d2;
#10 word33='d0;#10 word34='d2;
#10 word34='d0;#10 word35='d2;
#10 word35='d0;#10 word0='d4;
#10 word0='d0;#10 word1='d4;
#10 word1='d0;#10 word2='d4;
#10 word2='d0;#10 word3='d4;
#10 word3='d0;#10 word4='d4;
#10 word4='d0;#10 word5='d4;
#10 word5='d0;#10 word6='d4;
#10 word6='d0;#10 word7='d4;
#10 word7='d0;#10 word8='d4;
#10 word8='d0;#10 word9='d4;
#10 word9='d0;#10 word10='d4;
#10 word10='d0;#10 word11='d4;
#10 word11='d0;#10 word12='d4;
#10 word12='d0;#10 word13='d4;
#10 word13='d0;#10 word14='d4;
#10 word14='d0;#10 word15='d4;
#10 word15='d0;#10 word16='d4;
#10 word16='d0;#10 word17='d4;
#10 word17='d0;#10 word18='d4;
#10 word18='d0;#10 word19='d4;
#10 word19='d0;#10 word20='d4;
#10 word20='d0;#10 word21='d4;
#10 word21='d0;#10 word22='d4;
#10 word22='d0;#10 word23='d4;
#10 word23='d0;#10 word24='d4;
#10 word24='d0;#10 word25='d4;
#10 word25='d0;#10 word26='d4;
#10 word26='d0;#10 word27='d4;
#10 word27='d0;#10 word28='d4;
#10 word28='d0;#10 word29='d4;
#10 word29='d0;#10 word30='d4;
#10 word30='d0;#10 word31='d4;
#10 word31='d0;#10 word32='d4;
#10 word32='d0;#10 word33='d4;
#10 word33='d0;#10 word34='d4;
#10 word34='d0;#10 word35='d4;
#10 word35='d0;#10 word0='d8;
#10 word0='d0;#10 word1='d8;
#10 word1='d0;#10 word2='d8;
#10 word2='d0;#10 word3='d8;
#10 word3='d0;#10 word4='d8;
#10 word4='d0;#10 word5='d8;
#10 word5='d0;#10 word6='d8;
#10 word6='d0;#10 word7='d8;
#10 word7='d0;#10 word8='d8;
#10 word8='d0;#10 word9='d8;
#10 word9='d0;#10 word10='d8;
#10 word10='d0;#10 word11='d8;
#10 word11='d0;#10 word12='d8;
#10 word12='d0;#10 word13='d8;
#10 word13='d0;#10 word14='d8;
#10 word14='d0;#10 word15='d8;
#10 word15='d0;#10 word16='d8;
#10 word16='d0;#10 word17='d8;
#10 word17='d0;#10 word18='d8;
#10 word18='d0;#10 word19='d8;
#10 word19='d0;#10 word20='d8;
#10 word20='d0;#10 word21='d8;
#10 word21='d0;#10 word22='d8;
#10 word22='d0;#10 word23='d8;
#10 word23='d0;#10 word24='d8;
#10 word24='d0;#10 word25='d8;
#10 word25='d0;#10 word26='d8;
#10 word26='d0;#10 word27='d8;
#10 word27='d0;#10 word28='d8;
#10 word28='d0;#10 word29='d8;
#10 word29='d0;#10 word30='d8;
#10 word30='d0;#10 word31='d8;
#10 word31='d0;#10 word32='d8;
#10 word32='d0;#10 word33='d8;
#10 word33='d0;#10 word34='d8;
#10 word34='d0;#10 word35='d8;
#10 word35='d0;#10 word0='d16;
#10 word0='d0;#10 word1='d16;
#10 word1='d0;#10 word2='d16;
#10 word2='d0;#10 word3='d16;
#10 word3='d0;#10 word4='d16;
#10 word4='d0;#10 word5='d16;
#10 word5='d0;#10 word6='d16;
#10 word6='d0;#10 word7='d16;
#10 word7='d0;#10 word8='d16;
#10 word8='d0;#10 word9='d16;
#10 word9='d0;#10 word10='d16;
#10 word10='d0;#10 word11='d16;
#10 word11='d0;#10 word12='d16;
#10 word12='d0;#10 word13='d16;
#10 word13='d0;#10 word14='d16;
#10 word14='d0;#10 word15='d16;
#10 word15='d0;#10 word16='d16;
#10 word16='d0;#10 word17='d16;
#10 word17='d0;#10 word18='d16;
#10 word18='d0;#10 word19='d16;
#10 word19='d0;#10 word20='d16;
#10 word20='d0;#10 word21='d16;
#10 word21='d0;#10 word22='d16;
#10 word22='d0;#10 word23='d16;
#10 word23='d0;#10 word24='d16;
#10 word24='d0;#10 word25='d16;
#10 word25='d0;#10 word26='d16;
#10 word26='d0;#10 word27='d16;
#10 word27='d0;#10 word28='d16;
#10 word28='d0;#10 word29='d16;
#10 word29='d0;#10 word30='d16;
#10 word30='d0;#10 word31='d16;
#10 word31='d0;#10 word32='d16;
#10 word32='d0;#10 word33='d16;
#10 word33='d0;#10 word34='d16;
#10 word34='d0;#10 word35='d16;
#10 word35='d0;#10 word0='d32;
#10 word0='d0;#10 word1='d32;
#10 word1='d0;#10 word2='d32;
#10 word2='d0;#10 word3='d32;
#10 word3='d0;#10 word4='d32;
#10 word4='d0;#10 word5='d32;
#10 word5='d0;#10 word6='d32;
#10 word6='d0;#10 word7='d32;
#10 word7='d0;#10 word8='d32;
#10 word8='d0;#10 word9='d32;
#10 word9='d0;#10 word10='d32;
#10 word10='d0;#10 word11='d32;
#10 word11='d0;#10 word12='d32;
#10 word12='d0;#10 word13='d32;
#10 word13='d0;#10 word14='d32;
#10 word14='d0;#10 word15='d32;
#10 word15='d0;#10 word16='d32;
#10 word16='d0;#10 word17='d32;
#10 word17='d0;#10 word18='d32;
#10 word18='d0;#10 word19='d32;
#10 word19='d0;#10 word20='d32;
#10 word20='d0;#10 word21='d32;
#10 word21='d0;#10 word22='d32;
#10 word22='d0;#10 word23='d32;
#10 word23='d0;#10 word24='d32;
#10 word24='d0;#10 word25='d32;
#10 word25='d0;#10 word26='d32;
#10 word26='d0;#10 word27='d32;
#10 word27='d0;#10 word28='d32;
#10 word28='d0;#10 word29='d32;
#10 word29='d0;#10 word30='d32;
#10 word30='d0;#10 word31='d32;
#10 word31='d0;#10 word32='d32;
#10 word32='d0;#10 word33='d32;
#10 word33='d0;#10 word34='d32;
#10 word34='d0;#10 word35='d32;
#10 word35='d0;#10 word0='d12;
#10 word0='d0;#10 word1='d12;
#10 word1='d0;#10 word2='d12;
#10 word2='d0;#10 word3='d12;
#10 word3='d0;#10 word4='d12;
#10 word4='d0;#10 word5='d12;
#10 word5='d0;#10 word6='d12;
#10 word6='d0;#10 word7='d12;
#10 word7='d0;#10 word8='d12;
#10 word8='d0;#10 word9='d12;
#10 word9='d0;#10 word10='d12;
#10 word10='d0;#10 word11='d12;
#10 word11='d0;#10 word12='d12;
#10 word12='d0;#10 word13='d12;
#10 word13='d0;#10 word14='d12;
#10 word14='d0;#10 word15='d12;
#10 word15='d0;#10 word16='d12;
#10 word16='d0;#10 word17='d12;
#10 word17='d0;#10 word18='d12;
#10 word18='d0;#10 word19='d12;
#10 word19='d0;#10 word20='d12;
#10 word20='d0;#10 word21='d12;
#10 word21='d0;#10 word22='d12;
#10 word22='d0;#10 word23='d12;
#10 word23='d0;#10 word24='d12;
#10 word24='d0;#10 word25='d12;
#10 word25='d0;#10 word26='d12;
#10 word26='d0;#10 word27='d12;
#10 word27='d0;#10 word28='d12;
#10 word28='d0;#10 word29='d12;
#10 word29='d0;#10 word30='d12;
#10 word30='d0;#10 word31='d12;
#10 word31='d0;#10 word32='d12;
#10 word32='d0;#10 word33='d12;
#10 word33='d0;#10 word34='d12;
#10 word34='d0;#10 word35='d12;
#10 word35='d0;#10 word0='d15;
#10 word0='d0;#10 word1='d15;
#10 word1='d0;#10 word2='d15;
#10 word2='d0;#10 word3='d15;
#10 word3='d0;#10 word4='d15;
#10 word4='d0;#10 word5='d15;
#10 word5='d0;#10 word6='d15;
#10 word6='d0;#10 word7='d15;
#10 word7='d0;#10 word8='d15;
#10 word8='d0;#10 word9='d15;
#10 word9='d0;#10 word10='d15;
#10 word10='d0;#10 word11='d15;
#10 word11='d0;#10 word12='d15;
#10 word12='d0;#10 word13='d15;
#10 word13='d0;#10 word14='d15;
#10 word14='d0;#10 word15='d15;
#10 word15='d0;#10 word16='d15;
#10 word16='d0;#10 word17='d15;
#10 word17='d0;#10 word18='d15;
#10 word18='d0;#10 word19='d15;
#10 word19='d0;#10 word20='d15;
#10 word20='d0;#10 word21='d15;
#10 word21='d0;#10 word22='d15;
#10 word22='d0;#10 word23='d15;
#10 word23='d0;#10 word24='d15;
#10 word24='d0;#10 word25='d15;
#10 word25='d0;#10 word26='d15;
#10 word26='d0;#10 word27='d15;
#10 word27='d0;#10 word28='d15;
#10 word28='d0;#10 word29='d15;
#10 word29='d0;#10 word30='d15;
#10 word30='d0;#10 word31='d15;
#10 word31='d0;#10 word32='d15;
#10 word32='d0;#10 word33='d15;
#10 word33='d0;#10 word34='d15;
#10 word34='d0;#10 word35='d15;
#10 word35='d0;#10 word0='d9;
#10 word0='d0;#10 word1='d9;
#10 word1='d0;#10 word2='d9;
#10 word2='d0;#10 word3='d9;
#10 word3='d0;#10 word4='d9;
#10 word4='d0;#10 word5='d9;
#10 word5='d0;#10 word6='d9;
#10 word6='d0;#10 word7='d9;
#10 word7='d0;#10 word8='d9;
#10 word8='d0;#10 word9='d9;
#10 word9='d0;#10 word10='d9;
#10 word10='d0;#10 word11='d9;
#10 word11='d0;#10 word12='d9;
#10 word12='d0;#10 word13='d9;
#10 word13='d0;#10 word14='d9;
#10 word14='d0;#10 word15='d9;
#10 word15='d0;#10 word16='d9;
#10 word16='d0;#10 word17='d9;
#10 word17='d0;#10 word18='d9;
#10 word18='d0;#10 word19='d9;
#10 word19='d0;#10 word20='d9;
#10 word20='d0;#10 word21='d9;
#10 word21='d0;#10 word22='d9;
#10 word22='d0;#10 word23='d9;
#10 word23='d0;#10 word24='d9;
#10 word24='d0;#10 word25='d9;
#10 word25='d0;#10 word26='d9;
#10 word26='d0;#10 word27='d9;
#10 word27='d0;#10 word28='d9;
#10 word28='d0;#10 word29='d9;
#10 word29='d0;#10 word30='d9;
#10 word30='d0;#10 word31='d9;
#10 word31='d0;#10 word32='d9;
#10 word32='d0;#10 word33='d9;
#10 word33='d0;#10 word34='d9;
#10 word34='d0;#10 word35='d9;
#10 word35='d0;#10 word0='d5;
#10 word0='d0;#10 word1='d5;
#10 word1='d0;#10 word2='d5;
#10 word2='d0;#10 word3='d5;
#10 word3='d0;#10 word4='d5;
#10 word4='d0;#10 word5='d5;
#10 word5='d0;#10 word6='d5;
#10 word6='d0;#10 word7='d5;
#10 word7='d0;#10 word8='d5;
#10 word8='d0;#10 word9='d5;
#10 word9='d0;#10 word10='d5;
#10 word10='d0;#10 word11='d5;
#10 word11='d0;#10 word12='d5;
#10 word12='d0;#10 word13='d5;
#10 word13='d0;#10 word14='d5;
#10 word14='d0;#10 word15='d5;
#10 word15='d0;#10 word16='d5;
#10 word16='d0;#10 word17='d5;
#10 word17='d0;#10 word18='d5;
#10 word18='d0;#10 word19='d5;
#10 word19='d0;#10 word20='d5;
#10 word20='d0;#10 word21='d5;
#10 word21='d0;#10 word22='d5;
#10 word22='d0;#10 word23='d5;
#10 word23='d0;#10 word24='d5;
#10 word24='d0;#10 word25='d5;
#10 word25='d0;#10 word26='d5;
#10 word26='d0;#10 word27='d5;
#10 word27='d0;#10 word28='d5;
#10 word28='d0;#10 word29='d5;
#10 word29='d0;#10 word30='d5;
#10 word30='d0;#10 word31='d5;
#10 word31='d0;#10 word32='d5;
#10 word32='d0;#10 word33='d5;
#10 word33='d0;#10 word34='d5;
#10 word34='d0;#10 word35='d5;
#10 word35='d0;#10 word0='d29;
#10 word0='d0;#10 word1='d29;
#10 word1='d0;#10 word2='d29;
#10 word2='d0;#10 word3='d29;
#10 word3='d0;#10 word4='d29;
#10 word4='d0;#10 word5='d29;
#10 word5='d0;#10 word6='d29;
#10 word6='d0;#10 word7='d29;
#10 word7='d0;#10 word8='d29;
#10 word8='d0;#10 word9='d29;
#10 word9='d0;#10 word10='d29;
#10 word10='d0;#10 word11='d29;
#10 word11='d0;#10 word12='d29;
#10 word12='d0;#10 word13='d29;
#10 word13='d0;#10 word14='d29;
#10 word14='d0;#10 word15='d29;
#10 word15='d0;#10 word16='d29;
#10 word16='d0;#10 word17='d29;
#10 word17='d0;#10 word18='d29;
#10 word18='d0;#10 word19='d29;
#10 word19='d0;#10 word20='d29;
#10 word20='d0;#10 word21='d29;
#10 word21='d0;#10 word22='d29;
#10 word22='d0;#10 word23='d29;
#10 word23='d0;#10 word24='d29;
#10 word24='d0;#10 word25='d29;
#10 word25='d0;#10 word26='d29;
#10 word26='d0;#10 word27='d29;
#10 word27='d0;#10 word28='d29;
#10 word28='d0;#10 word29='d29;
#10 word29='d0;#10 word30='d29;
#10 word30='d0;#10 word31='d29;
#10 word31='d0;#10 word32='d29;
#10 word32='d0;#10 word33='d29;
#10 word33='d0;#10 word34='d29;
#10 word34='d0;#10 word35='d29;
#10 word35='d0;#10 word0='d45;
#10 word0='d0;#10 word1='d45;
#10 word1='d0;#10 word2='d45;
#10 word2='d0;#10 word3='d45;
#10 word3='d0;#10 word4='d45;
#10 word4='d0;#10 word5='d45;
#10 word5='d0;#10 word6='d45;
#10 word6='d0;#10 word7='d45;
#10 word7='d0;#10 word8='d45;
#10 word8='d0;#10 word9='d45;
#10 word9='d0;#10 word10='d45;
#10 word10='d0;#10 word11='d45;
#10 word11='d0;#10 word12='d45;
#10 word12='d0;#10 word13='d45;
#10 word13='d0;#10 word14='d45;
#10 word14='d0;#10 word15='d45;
#10 word15='d0;#10 word16='d45;
#10 word16='d0;#10 word17='d45;
#10 word17='d0;#10 word18='d45;
#10 word18='d0;#10 word19='d45;
#10 word19='d0;#10 word20='d45;
#10 word20='d0;#10 word21='d45;
#10 word21='d0;#10 word22='d45;
#10 word22='d0;#10 word23='d45;
#10 word23='d0;#10 word24='d45;
#10 word24='d0;#10 word25='d45;
#10 word25='d0;#10 word26='d45;
#10 word26='d0;#10 word27='d45;
#10 word27='d0;#10 word28='d45;
#10 word28='d0;#10 word29='d45;
#10 word29='d0;#10 word30='d45;
#10 word30='d0;#10 word31='d45;
#10 word31='d0;#10 word32='d45;
#10 word32='d0;#10 word33='d45;
#10 word33='d0;#10 word34='d45;
#10 word34='d0;#10 word35='d45;
#10 word35='d0;#10 word0='d27;
#10 word0='d0;#10 word1='d27;
#10 word1='d0;#10 word2='d27;
#10 word2='d0;#10 word3='d27;
#10 word3='d0;#10 word4='d27;
#10 word4='d0;#10 word5='d27;
#10 word5='d0;#10 word6='d27;
#10 word6='d0;#10 word7='d27;
#10 word7='d0;#10 word8='d27;
#10 word8='d0;#10 word9='d27;
#10 word9='d0;#10 word10='d27;
#10 word10='d0;#10 word11='d27;
#10 word11='d0;#10 word12='d27;
#10 word12='d0;#10 word13='d27;
#10 word13='d0;#10 word14='d27;
#10 word14='d0;#10 word15='d27;
#10 word15='d0;#10 word16='d27;
#10 word16='d0;#10 word17='d27;
#10 word17='d0;#10 word18='d27;
#10 word18='d0;#10 word19='d27;
#10 word19='d0;#10 word20='d27;
#10 word20='d0;#10 word21='d27;
#10 word21='d0;#10 word22='d27;
#10 word22='d0;#10 word23='d27;
#10 word23='d0;#10 word24='d27;
#10 word24='d0;#10 word25='d27;
#10 word25='d0;#10 word26='d27;
#10 word26='d0;#10 word27='d27;
#10 word27='d0;#10 word28='d27;
#10 word28='d0;#10 word29='d27;
#10 word29='d0;#10 word30='d27;
#10 word30='d0;#10 word31='d27;
#10 word31='d0;#10 word32='d27;
#10 word32='d0;#10 word33='d27;
#10 word33='d0;#10 word34='d27;
#10 word34='d0;#10 word35='d27;
#10 word35='d0;#10 word0='d24;
#10 word0='d0;#10 word1='d24;
#10 word1='d0;#10 word2='d24;
#10 word2='d0;#10 word3='d24;
#10 word3='d0;#10 word4='d24;
#10 word4='d0;#10 word5='d24;
#10 word5='d0;#10 word6='d24;
#10 word6='d0;#10 word7='d24;
#10 word7='d0;#10 word8='d24;
#10 word8='d0;#10 word9='d24;
#10 word9='d0;#10 word10='d24;
#10 word10='d0;#10 word11='d24;
#10 word11='d0;#10 word12='d24;
#10 word12='d0;#10 word13='d24;
#10 word13='d0;#10 word14='d24;
#10 word14='d0;#10 word15='d24;
#10 word15='d0;#10 word16='d24;
#10 word16='d0;#10 word17='d24;
#10 word17='d0;#10 word18='d24;
#10 word18='d0;#10 word19='d24;
#10 word19='d0;#10 word20='d24;
#10 word20='d0;#10 word21='d24;
#10 word21='d0;#10 word22='d24;
#10 word22='d0;#10 word23='d24;
#10 word23='d0;#10 word24='d24;
#10 word24='d0;#10 word25='d24;
#10 word25='d0;#10 word26='d24;
#10 word26='d0;#10 word27='d24;
#10 word27='d0;#10 word28='d24;
#10 word28='d0;#10 word29='d24;
#10 word29='d0;#10 word30='d24;
#10 word30='d0;#10 word31='d24;
#10 word31='d0;#10 word32='d24;
#10 word32='d0;#10 word33='d24;
#10 word33='d0;#10 word34='d24;
#10 word34='d0;#10 word35='d24;
#10 word35='d0;#10 word0='d30;
#10 word0='d0;#10 word1='d30;
#10 word1='d0;#10 word2='d30;
#10 word2='d0;#10 word3='d30;
#10 word3='d0;#10 word4='d30;
#10 word4='d0;#10 word5='d30;
#10 word5='d0;#10 word6='d30;
#10 word6='d0;#10 word7='d30;
#10 word7='d0;#10 word8='d30;
#10 word8='d0;#10 word9='d30;
#10 word9='d0;#10 word10='d30;
#10 word10='d0;#10 word11='d30;
#10 word11='d0;#10 word12='d30;
#10 word12='d0;#10 word13='d30;
#10 word13='d0;#10 word14='d30;
#10 word14='d0;#10 word15='d30;
#10 word15='d0;#10 word16='d30;
#10 word16='d0;#10 word17='d30;
#10 word17='d0;#10 word18='d30;
#10 word18='d0;#10 word19='d30;
#10 word19='d0;#10 word20='d30;
#10 word20='d0;#10 word21='d30;
#10 word21='d0;#10 word22='d30;
#10 word22='d0;#10 word23='d30;
#10 word23='d0;#10 word24='d30;
#10 word24='d0;#10 word25='d30;
#10 word25='d0;#10 word26='d30;
#10 word26='d0;#10 word27='d30;
#10 word27='d0;#10 word28='d30;
#10 word28='d0;#10 word29='d30;
#10 word29='d0;#10 word30='d30;
#10 word30='d0;#10 word31='d30;
#10 word31='d0;#10 word32='d30;
#10 word32='d0;#10 word33='d30;
#10 word33='d0;#10 word34='d30;
#10 word34='d0;#10 word35='d30;
#10 word35='d0;#10 word0='d18;
#10 word0='d0;#10 word1='d18;
#10 word1='d0;#10 word2='d18;
#10 word2='d0;#10 word3='d18;
#10 word3='d0;#10 word4='d18;
#10 word4='d0;#10 word5='d18;
#10 word5='d0;#10 word6='d18;
#10 word6='d0;#10 word7='d18;
#10 word7='d0;#10 word8='d18;
#10 word8='d0;#10 word9='d18;
#10 word9='d0;#10 word10='d18;
#10 word10='d0;#10 word11='d18;
#10 word11='d0;#10 word12='d18;
#10 word12='d0;#10 word13='d18;
#10 word13='d0;#10 word14='d18;
#10 word14='d0;#10 word15='d18;
#10 word15='d0;#10 word16='d18;
#10 word16='d0;#10 word17='d18;
#10 word17='d0;#10 word18='d18;
#10 word18='d0;#10 word19='d18;
#10 word19='d0;#10 word20='d18;
#10 word20='d0;#10 word21='d18;
#10 word21='d0;#10 word22='d18;
#10 word22='d0;#10 word23='d18;
#10 word23='d0;#10 word24='d18;
#10 word24='d0;#10 word25='d18;
#10 word25='d0;#10 word26='d18;
#10 word26='d0;#10 word27='d18;
#10 word27='d0;#10 word28='d18;
#10 word28='d0;#10 word29='d18;
#10 word29='d0;#10 word30='d18;
#10 word30='d0;#10 word31='d18;
#10 word31='d0;#10 word32='d18;
#10 word32='d0;#10 word33='d18;
#10 word33='d0;#10 word34='d18;
#10 word34='d0;#10 word35='d18;
#10 word35='d0;#10 word0='d10;
#10 word0='d0;#10 word1='d10;
#10 word1='d0;#10 word2='d10;
#10 word2='d0;#10 word3='d10;
#10 word3='d0;#10 word4='d10;
#10 word4='d0;#10 word5='d10;
#10 word5='d0;#10 word6='d10;
#10 word6='d0;#10 word7='d10;
#10 word7='d0;#10 word8='d10;
#10 word8='d0;#10 word9='d10;
#10 word9='d0;#10 word10='d10;
#10 word10='d0;#10 word11='d10;
#10 word11='d0;#10 word12='d10;
#10 word12='d0;#10 word13='d10;
#10 word13='d0;#10 word14='d10;
#10 word14='d0;#10 word15='d10;
#10 word15='d0;#10 word16='d10;
#10 word16='d0;#10 word17='d10;
#10 word17='d0;#10 word18='d10;
#10 word18='d0;#10 word19='d10;
#10 word19='d0;#10 word20='d10;
#10 word20='d0;#10 word21='d10;
#10 word21='d0;#10 word22='d10;
#10 word22='d0;#10 word23='d10;
#10 word23='d0;#10 word24='d10;
#10 word24='d0;#10 word25='d10;
#10 word25='d0;#10 word26='d10;
#10 word26='d0;#10 word27='d10;
#10 word27='d0;#10 word28='d10;
#10 word28='d0;#10 word29='d10;
#10 word29='d0;#10 word30='d10;
#10 word30='d0;#10 word31='d10;
#10 word31='d0;#10 word32='d10;
#10 word32='d0;#10 word33='d10;
#10 word33='d0;#10 word34='d10;
#10 word34='d0;#10 word35='d10;
#10 word35='d0;#10 word0='d58;
#10 word0='d0;#10 word1='d58;
#10 word1='d0;#10 word2='d58;
#10 word2='d0;#10 word3='d58;
#10 word3='d0;#10 word4='d58;
#10 word4='d0;#10 word5='d58;
#10 word5='d0;#10 word6='d58;
#10 word6='d0;#10 word7='d58;
#10 word7='d0;#10 word8='d58;
#10 word8='d0;#10 word9='d58;
#10 word9='d0;#10 word10='d58;
#10 word10='d0;#10 word11='d58;
#10 word11='d0;#10 word12='d58;
#10 word12='d0;#10 word13='d58;
#10 word13='d0;#10 word14='d58;
#10 word14='d0;#10 word15='d58;
#10 word15='d0;#10 word16='d58;
#10 word16='d0;#10 word17='d58;
#10 word17='d0;#10 word18='d58;
#10 word18='d0;#10 word19='d58;
#10 word19='d0;#10 word20='d58;
#10 word20='d0;#10 word21='d58;
#10 word21='d0;#10 word22='d58;
#10 word22='d0;#10 word23='d58;
#10 word23='d0;#10 word24='d58;
#10 word24='d0;#10 word25='d58;
#10 word25='d0;#10 word26='d58;
#10 word26='d0;#10 word27='d58;
#10 word27='d0;#10 word28='d58;
#10 word28='d0;#10 word29='d58;
#10 word29='d0;#10 word30='d58;
#10 word30='d0;#10 word31='d58;
#10 word31='d0;#10 word32='d58;
#10 word32='d0;#10 word33='d58;
#10 word33='d0;#10 word34='d58;
#10 word34='d0;#10 word35='d58;
#10 word35='d0;#10 word0='d38;
#10 word0='d0;#10 word1='d38;
#10 word1='d0;#10 word2='d38;
#10 word2='d0;#10 word3='d38;
#10 word3='d0;#10 word4='d38;
#10 word4='d0;#10 word5='d38;
#10 word5='d0;#10 word6='d38;
#10 word6='d0;#10 word7='d38;
#10 word7='d0;#10 word8='d38;
#10 word8='d0;#10 word9='d38;
#10 word9='d0;#10 word10='d38;
#10 word10='d0;#10 word11='d38;
#10 word11='d0;#10 word12='d38;
#10 word12='d0;#10 word13='d38;
#10 word13='d0;#10 word14='d38;
#10 word14='d0;#10 word15='d38;
#10 word15='d0;#10 word16='d38;
#10 word16='d0;#10 word17='d38;
#10 word17='d0;#10 word18='d38;
#10 word18='d0;#10 word19='d38;
#10 word19='d0;#10 word20='d38;
#10 word20='d0;#10 word21='d38;
#10 word21='d0;#10 word22='d38;
#10 word22='d0;#10 word23='d38;
#10 word23='d0;#10 word24='d38;
#10 word24='d0;#10 word25='d38;
#10 word25='d0;#10 word26='d38;
#10 word26='d0;#10 word27='d38;
#10 word27='d0;#10 word28='d38;
#10 word28='d0;#10 word29='d38;
#10 word29='d0;#10 word30='d38;
#10 word30='d0;#10 word31='d38;
#10 word31='d0;#10 word32='d38;
#10 word32='d0;#10 word33='d38;
#10 word33='d0;#10 word34='d38;
#10 word34='d0;#10 word35='d38;
#10 word35='d0;#10 word0='d37;
#10 word0='d0;#10 word1='d37;
#10 word1='d0;#10 word2='d37;
#10 word2='d0;#10 word3='d37;
#10 word3='d0;#10 word4='d37;
#10 word4='d0;#10 word5='d37;
#10 word5='d0;#10 word6='d37;
#10 word6='d0;#10 word7='d37;
#10 word7='d0;#10 word8='d37;
#10 word8='d0;#10 word9='d37;
#10 word9='d0;#10 word10='d37;
#10 word10='d0;#10 word11='d37;
#10 word11='d0;#10 word12='d37;
#10 word12='d0;#10 word13='d37;
#10 word13='d0;#10 word14='d37;
#10 word14='d0;#10 word15='d37;
#10 word15='d0;#10 word16='d37;
#10 word16='d0;#10 word17='d37;
#10 word17='d0;#10 word18='d37;
#10 word18='d0;#10 word19='d37;
#10 word19='d0;#10 word20='d37;
#10 word20='d0;#10 word21='d37;
#10 word21='d0;#10 word22='d37;
#10 word22='d0;#10 word23='d37;
#10 word23='d0;#10 word24='d37;
#10 word24='d0;#10 word25='d37;
#10 word25='d0;#10 word26='d37;
#10 word26='d0;#10 word27='d37;
#10 word27='d0;#10 word28='d37;
#10 word28='d0;#10 word29='d37;
#10 word29='d0;#10 word30='d37;
#10 word30='d0;#10 word31='d37;
#10 word31='d0;#10 word32='d37;
#10 word32='d0;#10 word33='d37;
#10 word33='d0;#10 word34='d37;
#10 word34='d0;#10 word35='d37;
#10 word35='d0;#10 word0='d35;
#10 word0='d0;#10 word1='d35;
#10 word1='d0;#10 word2='d35;
#10 word2='d0;#10 word3='d35;
#10 word3='d0;#10 word4='d35;
#10 word4='d0;#10 word5='d35;
#10 word5='d0;#10 word6='d35;
#10 word6='d0;#10 word7='d35;
#10 word7='d0;#10 word8='d35;
#10 word8='d0;#10 word9='d35;
#10 word9='d0;#10 word10='d35;
#10 word10='d0;#10 word11='d35;
#10 word11='d0;#10 word12='d35;
#10 word12='d0;#10 word13='d35;
#10 word13='d0;#10 word14='d35;
#10 word14='d0;#10 word15='d35;
#10 word15='d0;#10 word16='d35;
#10 word16='d0;#10 word17='d35;
#10 word17='d0;#10 word18='d35;
#10 word18='d0;#10 word19='d35;
#10 word19='d0;#10 word20='d35;
#10 word20='d0;#10 word21='d35;
#10 word21='d0;#10 word22='d35;
#10 word22='d0;#10 word23='d35;
#10 word23='d0;#10 word24='d35;
#10 word24='d0;#10 word25='d35;
#10 word25='d0;#10 word26='d35;
#10 word26='d0;#10 word27='d35;
#10 word27='d0;#10 word28='d35;
#10 word28='d0;#10 word29='d35;
#10 word29='d0;#10 word30='d35;
#10 word30='d0;#10 word31='d35;
#10 word31='d0;#10 word32='d35;
#10 word32='d0;#10 word33='d35;
#10 word33='d0;#10 word34='d35;
#10 word34='d0;#10 word35='d35;
#10 word35='d0;#10 word0='d47;
#10 word0='d0;#10 word1='d47;
#10 word1='d0;#10 word2='d47;
#10 word2='d0;#10 word3='d47;
#10 word3='d0;#10 word4='d47;
#10 word4='d0;#10 word5='d47;
#10 word5='d0;#10 word6='d47;
#10 word6='d0;#10 word7='d47;
#10 word7='d0;#10 word8='d47;
#10 word8='d0;#10 word9='d47;
#10 word9='d0;#10 word10='d47;
#10 word10='d0;#10 word11='d47;
#10 word11='d0;#10 word12='d47;
#10 word12='d0;#10 word13='d47;
#10 word13='d0;#10 word14='d47;
#10 word14='d0;#10 word15='d47;
#10 word15='d0;#10 word16='d47;
#10 word16='d0;#10 word17='d47;
#10 word17='d0;#10 word18='d47;
#10 word18='d0;#10 word19='d47;
#10 word19='d0;#10 word20='d47;
#10 word20='d0;#10 word21='d47;
#10 word21='d0;#10 word22='d47;
#10 word22='d0;#10 word23='d47;
#10 word23='d0;#10 word24='d47;
#10 word24='d0;#10 word25='d47;
#10 word25='d0;#10 word26='d47;
#10 word26='d0;#10 word27='d47;
#10 word27='d0;#10 word28='d47;
#10 word28='d0;#10 word29='d47;
#10 word29='d0;#10 word30='d47;
#10 word30='d0;#10 word31='d47;
#10 word31='d0;#10 word32='d47;
#10 word32='d0;#10 word33='d47;
#10 word33='d0;#10 word34='d47;
#10 word34='d0;#10 word35='d47;
#10 word35='d0;#10 word0='d55;
#10 word0='d0;#10 word1='d55;
#10 word1='d0;#10 word2='d55;
#10 word2='d0;#10 word3='d55;
#10 word3='d0;#10 word4='d55;
#10 word4='d0;#10 word5='d55;
#10 word5='d0;#10 word6='d55;
#10 word6='d0;#10 word7='d55;
#10 word7='d0;#10 word8='d55;
#10 word8='d0;#10 word9='d55;
#10 word9='d0;#10 word10='d55;
#10 word10='d0;#10 word11='d55;
#10 word11='d0;#10 word12='d55;
#10 word12='d0;#10 word13='d55;
#10 word13='d0;#10 word14='d55;
#10 word14='d0;#10 word15='d55;
#10 word15='d0;#10 word16='d55;
#10 word16='d0;#10 word17='d55;
#10 word17='d0;#10 word18='d55;
#10 word18='d0;#10 word19='d55;
#10 word19='d0;#10 word20='d55;
#10 word20='d0;#10 word21='d55;
#10 word21='d0;#10 word22='d55;
#10 word22='d0;#10 word23='d55;
#10 word23='d0;#10 word24='d55;
#10 word24='d0;#10 word25='d55;
#10 word25='d0;#10 word26='d55;
#10 word26='d0;#10 word27='d55;
#10 word27='d0;#10 word28='d55;
#10 word28='d0;#10 word29='d55;
#10 word29='d0;#10 word30='d55;
#10 word30='d0;#10 word31='d55;
#10 word31='d0;#10 word32='d55;
#10 word32='d0;#10 word33='d55;
#10 word33='d0;#10 word34='d55;
#10 word34='d0;#10 word35='d55;
#10 word35='d0;#10 word0='d7;
#10 word0='d0;#10 word1='d7;
#10 word1='d0;#10 word2='d7;
#10 word2='d0;#10 word3='d7;
#10 word3='d0;#10 word4='d7;
#10 word4='d0;#10 word5='d7;
#10 word5='d0;#10 word6='d7;
#10 word6='d0;#10 word7='d7;
#10 word7='d0;#10 word8='d7;
#10 word8='d0;#10 word9='d7;
#10 word9='d0;#10 word10='d7;
#10 word10='d0;#10 word11='d7;
#10 word11='d0;#10 word12='d7;
#10 word12='d0;#10 word13='d7;
#10 word13='d0;#10 word14='d7;
#10 word14='d0;#10 word15='d7;
#10 word15='d0;#10 word16='d7;
#10 word16='d0;#10 word17='d7;
#10 word17='d0;#10 word18='d7;
#10 word18='d0;#10 word19='d7;
#10 word19='d0;#10 word20='d7;
#10 word20='d0;#10 word21='d7;
#10 word21='d0;#10 word22='d7;
#10 word22='d0;#10 word23='d7;
#10 word23='d0;#10 word24='d7;
#10 word24='d0;#10 word25='d7;
#10 word25='d0;#10 word26='d7;
#10 word26='d0;#10 word27='d7;
#10 word27='d0;#10 word28='d7;
#10 word28='d0;#10 word29='d7;
#10 word29='d0;#10 word30='d7;
#10 word30='d0;#10 word31='d7;
#10 word31='d0;#10 word32='d7;
#10 word32='d0;#10 word33='d7;
#10 word33='d0;#10 word34='d7;
#10 word34='d0;#10 word35='d7;
#10 word35='d0;#10 word0='d53;
#10 word0='d0;#10 word1='d53;
#10 word1='d0;#10 word2='d53;
#10 word2='d0;#10 word3='d53;
#10 word3='d0;#10 word4='d53;
#10 word4='d0;#10 word5='d53;
#10 word5='d0;#10 word6='d53;
#10 word6='d0;#10 word7='d53;
#10 word7='d0;#10 word8='d53;
#10 word8='d0;#10 word9='d53;
#10 word9='d0;#10 word10='d53;
#10 word10='d0;#10 word11='d53;
#10 word11='d0;#10 word12='d53;
#10 word12='d0;#10 word13='d53;
#10 word13='d0;#10 word14='d53;
#10 word14='d0;#10 word15='d53;
#10 word15='d0;#10 word16='d53;
#10 word16='d0;#10 word17='d53;
#10 word17='d0;#10 word18='d53;
#10 word18='d0;#10 word19='d53;
#10 word19='d0;#10 word20='d53;
#10 word20='d0;#10 word21='d53;
#10 word21='d0;#10 word22='d53;
#10 word22='d0;#10 word23='d53;
#10 word23='d0;#10 word24='d53;
#10 word24='d0;#10 word25='d53;
#10 word25='d0;#10 word26='d53;
#10 word26='d0;#10 word27='d53;
#10 word27='d0;#10 word28='d53;
#10 word28='d0;#10 word29='d53;
#10 word29='d0;#10 word30='d53;
#10 word30='d0;#10 word31='d53;
#10 word31='d0;#10 word32='d53;
#10 word32='d0;#10 word33='d53;
#10 word33='d0;#10 word34='d53;
#10 word34='d0;#10 word35='d53;
#10 word35='d0;#10 word0='d54;
#10 word0='d0;#10 word1='d54;
#10 word1='d0;#10 word2='d54;
#10 word2='d0;#10 word3='d54;
#10 word3='d0;#10 word4='d54;
#10 word4='d0;#10 word5='d54;
#10 word5='d0;#10 word6='d54;
#10 word6='d0;#10 word7='d54;
#10 word7='d0;#10 word8='d54;
#10 word8='d0;#10 word9='d54;
#10 word9='d0;#10 word10='d54;
#10 word10='d0;#10 word11='d54;
#10 word11='d0;#10 word12='d54;
#10 word12='d0;#10 word13='d54;
#10 word13='d0;#10 word14='d54;
#10 word14='d0;#10 word15='d54;
#10 word15='d0;#10 word16='d54;
#10 word16='d0;#10 word17='d54;
#10 word17='d0;#10 word18='d54;
#10 word18='d0;#10 word19='d54;
#10 word19='d0;#10 word20='d54;
#10 word20='d0;#10 word21='d54;
#10 word21='d0;#10 word22='d54;
#10 word22='d0;#10 word23='d54;
#10 word23='d0;#10 word24='d54;
#10 word24='d0;#10 word25='d54;
#10 word25='d0;#10 word26='d54;
#10 word26='d0;#10 word27='d54;
#10 word27='d0;#10 word28='d54;
#10 word28='d0;#10 word29='d54;
#10 word29='d0;#10 word30='d54;
#10 word30='d0;#10 word31='d54;
#10 word31='d0;#10 word32='d54;
#10 word32='d0;#10 word33='d54;
#10 word33='d0;#10 word34='d54;
#10 word34='d0;#10 word35='d54;
#10 word35='d0;#10 word0='d48;
#10 word0='d0;#10 word1='d48;
#10 word1='d0;#10 word2='d48;
#10 word2='d0;#10 word3='d48;
#10 word3='d0;#10 word4='d48;
#10 word4='d0;#10 word5='d48;
#10 word5='d0;#10 word6='d48;
#10 word6='d0;#10 word7='d48;
#10 word7='d0;#10 word8='d48;
#10 word8='d0;#10 word9='d48;
#10 word9='d0;#10 word10='d48;
#10 word10='d0;#10 word11='d48;
#10 word11='d0;#10 word12='d48;
#10 word12='d0;#10 word13='d48;
#10 word13='d0;#10 word14='d48;
#10 word14='d0;#10 word15='d48;
#10 word15='d0;#10 word16='d48;
#10 word16='d0;#10 word17='d48;
#10 word17='d0;#10 word18='d48;
#10 word18='d0;#10 word19='d48;
#10 word19='d0;#10 word20='d48;
#10 word20='d0;#10 word21='d48;
#10 word21='d0;#10 word22='d48;
#10 word22='d0;#10 word23='d48;
#10 word23='d0;#10 word24='d48;
#10 word24='d0;#10 word25='d48;
#10 word25='d0;#10 word26='d48;
#10 word26='d0;#10 word27='d48;
#10 word27='d0;#10 word28='d48;
#10 word28='d0;#10 word29='d48;
#10 word29='d0;#10 word30='d48;
#10 word30='d0;#10 word31='d48;
#10 word31='d0;#10 word32='d48;
#10 word32='d0;#10 word33='d48;
#10 word33='d0;#10 word34='d48;
#10 word34='d0;#10 word35='d48;
#10 word35='d0;#10 word0='d60;
#10 word0='d0;#10 word1='d60;
#10 word1='d0;#10 word2='d60;
#10 word2='d0;#10 word3='d60;
#10 word3='d0;#10 word4='d60;
#10 word4='d0;#10 word5='d60;
#10 word5='d0;#10 word6='d60;
#10 word6='d0;#10 word7='d60;
#10 word7='d0;#10 word8='d60;
#10 word8='d0;#10 word9='d60;
#10 word9='d0;#10 word10='d60;
#10 word10='d0;#10 word11='d60;
#10 word11='d0;#10 word12='d60;
#10 word12='d0;#10 word13='d60;
#10 word13='d0;#10 word14='d60;
#10 word14='d0;#10 word15='d60;
#10 word15='d0;#10 word16='d60;
#10 word16='d0;#10 word17='d60;
#10 word17='d0;#10 word18='d60;
#10 word18='d0;#10 word19='d60;
#10 word19='d0;#10 word20='d60;
#10 word20='d0;#10 word21='d60;
#10 word21='d0;#10 word22='d60;
#10 word22='d0;#10 word23='d60;
#10 word23='d0;#10 word24='d60;
#10 word24='d0;#10 word25='d60;
#10 word25='d0;#10 word26='d60;
#10 word26='d0;#10 word27='d60;
#10 word27='d0;#10 word28='d60;
#10 word28='d0;#10 word29='d60;
#10 word29='d0;#10 word30='d60;
#10 word30='d0;#10 word31='d60;
#10 word31='d0;#10 word32='d60;
#10 word32='d0;#10 word33='d60;
#10 word33='d0;#10 word34='d60;
#10 word34='d0;#10 word35='d60;
#10 word35='d0;#10 word0='d36;
#10 word0='d0;#10 word1='d36;
#10 word1='d0;#10 word2='d36;
#10 word2='d0;#10 word3='d36;
#10 word3='d0;#10 word4='d36;
#10 word4='d0;#10 word5='d36;
#10 word5='d0;#10 word6='d36;
#10 word6='d0;#10 word7='d36;
#10 word7='d0;#10 word8='d36;
#10 word8='d0;#10 word9='d36;
#10 word9='d0;#10 word10='d36;
#10 word10='d0;#10 word11='d36;
#10 word11='d0;#10 word12='d36;
#10 word12='d0;#10 word13='d36;
#10 word13='d0;#10 word14='d36;
#10 word14='d0;#10 word15='d36;
#10 word15='d0;#10 word16='d36;
#10 word16='d0;#10 word17='d36;
#10 word17='d0;#10 word18='d36;
#10 word18='d0;#10 word19='d36;
#10 word19='d0;#10 word20='d36;
#10 word20='d0;#10 word21='d36;
#10 word21='d0;#10 word22='d36;
#10 word22='d0;#10 word23='d36;
#10 word23='d0;#10 word24='d36;
#10 word24='d0;#10 word25='d36;
#10 word25='d0;#10 word26='d36;
#10 word26='d0;#10 word27='d36;
#10 word27='d0;#10 word28='d36;
#10 word28='d0;#10 word29='d36;
#10 word29='d0;#10 word30='d36;
#10 word30='d0;#10 word31='d36;
#10 word31='d0;#10 word32='d36;
#10 word32='d0;#10 word33='d36;
#10 word33='d0;#10 word34='d36;
#10 word34='d0;#10 word35='d36;
#10 word35='d0;#10 word0='d20;
#10 word0='d0;#10 word1='d20;
#10 word1='d0;#10 word2='d20;
#10 word2='d0;#10 word3='d20;
#10 word3='d0;#10 word4='d20;
#10 word4='d0;#10 word5='d20;
#10 word5='d0;#10 word6='d20;
#10 word6='d0;#10 word7='d20;
#10 word7='d0;#10 word8='d20;
#10 word8='d0;#10 word9='d20;
#10 word9='d0;#10 word10='d20;
#10 word10='d0;#10 word11='d20;
#10 word11='d0;#10 word12='d20;
#10 word12='d0;#10 word13='d20;
#10 word13='d0;#10 word14='d20;
#10 word14='d0;#10 word15='d20;
#10 word15='d0;#10 word16='d20;
#10 word16='d0;#10 word17='d20;
#10 word17='d0;#10 word18='d20;
#10 word18='d0;#10 word19='d20;
#10 word19='d0;#10 word20='d20;
#10 word20='d0;#10 word21='d20;
#10 word21='d0;#10 word22='d20;
#10 word22='d0;#10 word23='d20;
#10 word23='d0;#10 word24='d20;
#10 word24='d0;#10 word25='d20;
#10 word25='d0;#10 word26='d20;
#10 word26='d0;#10 word27='d20;
#10 word27='d0;#10 word28='d20;
#10 word28='d0;#10 word29='d20;
#10 word29='d0;#10 word30='d20;
#10 word30='d0;#10 word31='d20;
#10 word31='d0;#10 word32='d20;
#10 word32='d0;#10 word33='d20;
#10 word33='d0;#10 word34='d20;
#10 word34='d0;#10 word35='d20;
#10 word35='d0;

    #20 $stop;
    end
endmodule
