module n19sys(input [8:0]IN0,input [8:0]IN1,output [4:0]OUT0,output [4:0]OUT1,