module convolution
    #(
        parameter   OUTPUT_BIT  =   19,
                    OUTPUT_NODE =   100,
                    DATA_WIDTH  =   19,
                    IMG_SZ    =   144
)
(
    input   clk,
    input   rst,
    input   [IMG_SZ*8-1:0]   img,
    input   valid,
    output  reg ready,
    output reg [OUTPUT_BIT*OUTPUT_NODE-1:0] layer_out
);

reg    signed [8-1:0]  in_buffer[0:IMG_SZ-1];
integer j;

always@(posedge clk)
    begin
        if(rst)
            begin
                for(j=0;j<IMG_SZ;j=j+1)
                    begin
                        in_buffer[j]<=0;
                    end
            end
        else
            begin
                for(j=0;j<IMG_SZ;j=j+1)
                    begin
                        in_buffer[j]<=img[j*8+:8];
                    end
            end
    end

//wire declatation
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight0;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight1;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight2;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight3;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight4;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight5;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight6;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight7;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight8;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight9;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight10;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight11;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight12;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight13;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight14;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight15;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight16;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight17;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight18;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight19;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight20;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight21;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight22;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight23;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight24;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight25;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight26;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight27;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight28;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight29;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight30;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight31;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight32;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight33;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight34;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight35;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight36;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight37;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight38;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight39;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight40;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight41;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight42;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight43;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight44;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight45;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight46;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight47;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight48;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight49;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight50;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight51;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight52;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight53;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight54;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight55;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight56;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight57;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight58;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight59;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight60;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight61;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight62;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight63;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight64;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight65;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight66;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight67;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight68;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight69;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight70;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight71;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight72;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight73;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight74;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight75;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight76;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight77;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight78;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight79;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight80;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight81;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight82;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight83;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight84;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight85;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight86;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight87;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight88;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight89;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight90;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight91;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight92;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight93;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight94;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight95;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight96;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight97;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight98;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight99;
assign in_buffer_weight0=$signed(in_buffer[0]*(41))+$signed(in_buffer[1]*(109))+$signed(in_buffer[2]*(108))+$signed(in_buffer[12]*(-58))+$signed(in_buffer[13]*(281))+$signed(in_buffer[14]*(143))+$signed(in_buffer[24]*(187))+$signed(in_buffer[25]*(188))+$signed(in_buffer[26]*(210));
assign in_buffer_weight1=$signed(in_buffer[1]*(41))+$signed(in_buffer[2]*(109))+$signed(in_buffer[3]*(108))+$signed(in_buffer[13]*(-58))+$signed(in_buffer[14]*(281))+$signed(in_buffer[15]*(143))+$signed(in_buffer[25]*(187))+$signed(in_buffer[26]*(188))+$signed(in_buffer[27]*(210));
assign in_buffer_weight2=$signed(in_buffer[2]*(41))+$signed(in_buffer[3]*(109))+$signed(in_buffer[4]*(108))+$signed(in_buffer[14]*(-58))+$signed(in_buffer[15]*(281))+$signed(in_buffer[16]*(143))+$signed(in_buffer[26]*(187))+$signed(in_buffer[27]*(188))+$signed(in_buffer[28]*(210));
assign in_buffer_weight3=$signed(in_buffer[3]*(41))+$signed(in_buffer[4]*(109))+$signed(in_buffer[5]*(108))+$signed(in_buffer[15]*(-58))+$signed(in_buffer[16]*(281))+$signed(in_buffer[17]*(143))+$signed(in_buffer[27]*(187))+$signed(in_buffer[28]*(188))+$signed(in_buffer[29]*(210));
assign in_buffer_weight4=$signed(in_buffer[4]*(41))+$signed(in_buffer[5]*(109))+$signed(in_buffer[6]*(108))+$signed(in_buffer[16]*(-58))+$signed(in_buffer[17]*(281))+$signed(in_buffer[18]*(143))+$signed(in_buffer[28]*(187))+$signed(in_buffer[29]*(188))+$signed(in_buffer[30]*(210));
assign in_buffer_weight5=$signed(in_buffer[5]*(41))+$signed(in_buffer[6]*(109))+$signed(in_buffer[7]*(108))+$signed(in_buffer[17]*(-58))+$signed(in_buffer[18]*(281))+$signed(in_buffer[19]*(143))+$signed(in_buffer[29]*(187))+$signed(in_buffer[30]*(188))+$signed(in_buffer[31]*(210));
assign in_buffer_weight6=$signed(in_buffer[6]*(41))+$signed(in_buffer[7]*(109))+$signed(in_buffer[8]*(108))+$signed(in_buffer[18]*(-58))+$signed(in_buffer[19]*(281))+$signed(in_buffer[20]*(143))+$signed(in_buffer[30]*(187))+$signed(in_buffer[31]*(188))+$signed(in_buffer[32]*(210));
assign in_buffer_weight7=$signed(in_buffer[7]*(41))+$signed(in_buffer[8]*(109))+$signed(in_buffer[9]*(108))+$signed(in_buffer[19]*(-58))+$signed(in_buffer[20]*(281))+$signed(in_buffer[21]*(143))+$signed(in_buffer[31]*(187))+$signed(in_buffer[32]*(188))+$signed(in_buffer[33]*(210));
assign in_buffer_weight8=$signed(in_buffer[8]*(41))+$signed(in_buffer[9]*(109))+$signed(in_buffer[10]*(108))+$signed(in_buffer[20]*(-58))+$signed(in_buffer[21]*(281))+$signed(in_buffer[22]*(143))+$signed(in_buffer[32]*(187))+$signed(in_buffer[33]*(188))+$signed(in_buffer[34]*(210));
assign in_buffer_weight9=$signed(in_buffer[9]*(41))+$signed(in_buffer[10]*(109))+$signed(in_buffer[11]*(108))+$signed(in_buffer[21]*(-58))+$signed(in_buffer[22]*(281))+$signed(in_buffer[23]*(143))+$signed(in_buffer[33]*(187))+$signed(in_buffer[34]*(188))+$signed(in_buffer[35]*(210));
assign in_buffer_weight10=$signed(in_buffer[12]*(41))+$signed(in_buffer[13]*(109))+$signed(in_buffer[14]*(108))+$signed(in_buffer[24]*(-58))+$signed(in_buffer[25]*(281))+$signed(in_buffer[26]*(143))+$signed(in_buffer[36]*(187))+$signed(in_buffer[37]*(188))+$signed(in_buffer[38]*(210));
assign in_buffer_weight11=$signed(in_buffer[13]*(41))+$signed(in_buffer[14]*(109))+$signed(in_buffer[15]*(108))+$signed(in_buffer[25]*(-58))+$signed(in_buffer[26]*(281))+$signed(in_buffer[27]*(143))+$signed(in_buffer[37]*(187))+$signed(in_buffer[38]*(188))+$signed(in_buffer[39]*(210));
assign in_buffer_weight12=$signed(in_buffer[14]*(41))+$signed(in_buffer[15]*(109))+$signed(in_buffer[16]*(108))+$signed(in_buffer[26]*(-58))+$signed(in_buffer[27]*(281))+$signed(in_buffer[28]*(143))+$signed(in_buffer[38]*(187))+$signed(in_buffer[39]*(188))+$signed(in_buffer[40]*(210));
assign in_buffer_weight13=$signed(in_buffer[15]*(41))+$signed(in_buffer[16]*(109))+$signed(in_buffer[17]*(108))+$signed(in_buffer[27]*(-58))+$signed(in_buffer[28]*(281))+$signed(in_buffer[29]*(143))+$signed(in_buffer[39]*(187))+$signed(in_buffer[40]*(188))+$signed(in_buffer[41]*(210));
assign in_buffer_weight14=$signed(in_buffer[16]*(41))+$signed(in_buffer[17]*(109))+$signed(in_buffer[18]*(108))+$signed(in_buffer[28]*(-58))+$signed(in_buffer[29]*(281))+$signed(in_buffer[30]*(143))+$signed(in_buffer[40]*(187))+$signed(in_buffer[41]*(188))+$signed(in_buffer[42]*(210));
assign in_buffer_weight15=$signed(in_buffer[17]*(41))+$signed(in_buffer[18]*(109))+$signed(in_buffer[19]*(108))+$signed(in_buffer[29]*(-58))+$signed(in_buffer[30]*(281))+$signed(in_buffer[31]*(143))+$signed(in_buffer[41]*(187))+$signed(in_buffer[42]*(188))+$signed(in_buffer[43]*(210));
assign in_buffer_weight16=$signed(in_buffer[18]*(41))+$signed(in_buffer[19]*(109))+$signed(in_buffer[20]*(108))+$signed(in_buffer[30]*(-58))+$signed(in_buffer[31]*(281))+$signed(in_buffer[32]*(143))+$signed(in_buffer[42]*(187))+$signed(in_buffer[43]*(188))+$signed(in_buffer[44]*(210));
assign in_buffer_weight17=$signed(in_buffer[19]*(41))+$signed(in_buffer[20]*(109))+$signed(in_buffer[21]*(108))+$signed(in_buffer[31]*(-58))+$signed(in_buffer[32]*(281))+$signed(in_buffer[33]*(143))+$signed(in_buffer[43]*(187))+$signed(in_buffer[44]*(188))+$signed(in_buffer[45]*(210));
assign in_buffer_weight18=$signed(in_buffer[20]*(41))+$signed(in_buffer[21]*(109))+$signed(in_buffer[22]*(108))+$signed(in_buffer[32]*(-58))+$signed(in_buffer[33]*(281))+$signed(in_buffer[34]*(143))+$signed(in_buffer[44]*(187))+$signed(in_buffer[45]*(188))+$signed(in_buffer[46]*(210));
assign in_buffer_weight19=$signed(in_buffer[21]*(41))+$signed(in_buffer[22]*(109))+$signed(in_buffer[23]*(108))+$signed(in_buffer[33]*(-58))+$signed(in_buffer[34]*(281))+$signed(in_buffer[35]*(143))+$signed(in_buffer[45]*(187))+$signed(in_buffer[46]*(188))+$signed(in_buffer[47]*(210));
assign in_buffer_weight20=$signed(in_buffer[24]*(41))+$signed(in_buffer[25]*(109))+$signed(in_buffer[26]*(108))+$signed(in_buffer[36]*(-58))+$signed(in_buffer[37]*(281))+$signed(in_buffer[38]*(143))+$signed(in_buffer[48]*(187))+$signed(in_buffer[49]*(188))+$signed(in_buffer[50]*(210));
assign in_buffer_weight21=$signed(in_buffer[25]*(41))+$signed(in_buffer[26]*(109))+$signed(in_buffer[27]*(108))+$signed(in_buffer[37]*(-58))+$signed(in_buffer[38]*(281))+$signed(in_buffer[39]*(143))+$signed(in_buffer[49]*(187))+$signed(in_buffer[50]*(188))+$signed(in_buffer[51]*(210));
assign in_buffer_weight22=$signed(in_buffer[26]*(41))+$signed(in_buffer[27]*(109))+$signed(in_buffer[28]*(108))+$signed(in_buffer[38]*(-58))+$signed(in_buffer[39]*(281))+$signed(in_buffer[40]*(143))+$signed(in_buffer[50]*(187))+$signed(in_buffer[51]*(188))+$signed(in_buffer[52]*(210));
assign in_buffer_weight23=$signed(in_buffer[27]*(41))+$signed(in_buffer[28]*(109))+$signed(in_buffer[29]*(108))+$signed(in_buffer[39]*(-58))+$signed(in_buffer[40]*(281))+$signed(in_buffer[41]*(143))+$signed(in_buffer[51]*(187))+$signed(in_buffer[52]*(188))+$signed(in_buffer[53]*(210));
assign in_buffer_weight24=$signed(in_buffer[28]*(41))+$signed(in_buffer[29]*(109))+$signed(in_buffer[30]*(108))+$signed(in_buffer[40]*(-58))+$signed(in_buffer[41]*(281))+$signed(in_buffer[42]*(143))+$signed(in_buffer[52]*(187))+$signed(in_buffer[53]*(188))+$signed(in_buffer[54]*(210));
assign in_buffer_weight25=$signed(in_buffer[29]*(41))+$signed(in_buffer[30]*(109))+$signed(in_buffer[31]*(108))+$signed(in_buffer[41]*(-58))+$signed(in_buffer[42]*(281))+$signed(in_buffer[43]*(143))+$signed(in_buffer[53]*(187))+$signed(in_buffer[54]*(188))+$signed(in_buffer[55]*(210));
assign in_buffer_weight26=$signed(in_buffer[30]*(41))+$signed(in_buffer[31]*(109))+$signed(in_buffer[32]*(108))+$signed(in_buffer[42]*(-58))+$signed(in_buffer[43]*(281))+$signed(in_buffer[44]*(143))+$signed(in_buffer[54]*(187))+$signed(in_buffer[55]*(188))+$signed(in_buffer[56]*(210));
assign in_buffer_weight27=$signed(in_buffer[31]*(41))+$signed(in_buffer[32]*(109))+$signed(in_buffer[33]*(108))+$signed(in_buffer[43]*(-58))+$signed(in_buffer[44]*(281))+$signed(in_buffer[45]*(143))+$signed(in_buffer[55]*(187))+$signed(in_buffer[56]*(188))+$signed(in_buffer[57]*(210));
assign in_buffer_weight28=$signed(in_buffer[32]*(41))+$signed(in_buffer[33]*(109))+$signed(in_buffer[34]*(108))+$signed(in_buffer[44]*(-58))+$signed(in_buffer[45]*(281))+$signed(in_buffer[46]*(143))+$signed(in_buffer[56]*(187))+$signed(in_buffer[57]*(188))+$signed(in_buffer[58]*(210));
assign in_buffer_weight29=$signed(in_buffer[33]*(41))+$signed(in_buffer[34]*(109))+$signed(in_buffer[35]*(108))+$signed(in_buffer[45]*(-58))+$signed(in_buffer[46]*(281))+$signed(in_buffer[47]*(143))+$signed(in_buffer[57]*(187))+$signed(in_buffer[58]*(188))+$signed(in_buffer[59]*(210));
assign in_buffer_weight30=$signed(in_buffer[36]*(41))+$signed(in_buffer[37]*(109))+$signed(in_buffer[38]*(108))+$signed(in_buffer[48]*(-58))+$signed(in_buffer[49]*(281))+$signed(in_buffer[50]*(143))+$signed(in_buffer[60]*(187))+$signed(in_buffer[61]*(188))+$signed(in_buffer[62]*(210));
assign in_buffer_weight31=$signed(in_buffer[37]*(41))+$signed(in_buffer[38]*(109))+$signed(in_buffer[39]*(108))+$signed(in_buffer[49]*(-58))+$signed(in_buffer[50]*(281))+$signed(in_buffer[51]*(143))+$signed(in_buffer[61]*(187))+$signed(in_buffer[62]*(188))+$signed(in_buffer[63]*(210));
assign in_buffer_weight32=$signed(in_buffer[38]*(41))+$signed(in_buffer[39]*(109))+$signed(in_buffer[40]*(108))+$signed(in_buffer[50]*(-58))+$signed(in_buffer[51]*(281))+$signed(in_buffer[52]*(143))+$signed(in_buffer[62]*(187))+$signed(in_buffer[63]*(188))+$signed(in_buffer[64]*(210));
assign in_buffer_weight33=$signed(in_buffer[39]*(41))+$signed(in_buffer[40]*(109))+$signed(in_buffer[41]*(108))+$signed(in_buffer[51]*(-58))+$signed(in_buffer[52]*(281))+$signed(in_buffer[53]*(143))+$signed(in_buffer[63]*(187))+$signed(in_buffer[64]*(188))+$signed(in_buffer[65]*(210));
assign in_buffer_weight34=$signed(in_buffer[40]*(41))+$signed(in_buffer[41]*(109))+$signed(in_buffer[42]*(108))+$signed(in_buffer[52]*(-58))+$signed(in_buffer[53]*(281))+$signed(in_buffer[54]*(143))+$signed(in_buffer[64]*(187))+$signed(in_buffer[65]*(188))+$signed(in_buffer[66]*(210));
assign in_buffer_weight35=$signed(in_buffer[41]*(41))+$signed(in_buffer[42]*(109))+$signed(in_buffer[43]*(108))+$signed(in_buffer[53]*(-58))+$signed(in_buffer[54]*(281))+$signed(in_buffer[55]*(143))+$signed(in_buffer[65]*(187))+$signed(in_buffer[66]*(188))+$signed(in_buffer[67]*(210));
assign in_buffer_weight36=$signed(in_buffer[42]*(41))+$signed(in_buffer[43]*(109))+$signed(in_buffer[44]*(108))+$signed(in_buffer[54]*(-58))+$signed(in_buffer[55]*(281))+$signed(in_buffer[56]*(143))+$signed(in_buffer[66]*(187))+$signed(in_buffer[67]*(188))+$signed(in_buffer[68]*(210));
assign in_buffer_weight37=$signed(in_buffer[43]*(41))+$signed(in_buffer[44]*(109))+$signed(in_buffer[45]*(108))+$signed(in_buffer[55]*(-58))+$signed(in_buffer[56]*(281))+$signed(in_buffer[57]*(143))+$signed(in_buffer[67]*(187))+$signed(in_buffer[68]*(188))+$signed(in_buffer[69]*(210));
assign in_buffer_weight38=$signed(in_buffer[44]*(41))+$signed(in_buffer[45]*(109))+$signed(in_buffer[46]*(108))+$signed(in_buffer[56]*(-58))+$signed(in_buffer[57]*(281))+$signed(in_buffer[58]*(143))+$signed(in_buffer[68]*(187))+$signed(in_buffer[69]*(188))+$signed(in_buffer[70]*(210));
assign in_buffer_weight39=$signed(in_buffer[45]*(41))+$signed(in_buffer[46]*(109))+$signed(in_buffer[47]*(108))+$signed(in_buffer[57]*(-58))+$signed(in_buffer[58]*(281))+$signed(in_buffer[59]*(143))+$signed(in_buffer[69]*(187))+$signed(in_buffer[70]*(188))+$signed(in_buffer[71]*(210));
assign in_buffer_weight40=$signed(in_buffer[48]*(41))+$signed(in_buffer[49]*(109))+$signed(in_buffer[50]*(108))+$signed(in_buffer[60]*(-58))+$signed(in_buffer[61]*(281))+$signed(in_buffer[62]*(143))+$signed(in_buffer[72]*(187))+$signed(in_buffer[73]*(188))+$signed(in_buffer[74]*(210));
assign in_buffer_weight41=$signed(in_buffer[49]*(41))+$signed(in_buffer[50]*(109))+$signed(in_buffer[51]*(108))+$signed(in_buffer[61]*(-58))+$signed(in_buffer[62]*(281))+$signed(in_buffer[63]*(143))+$signed(in_buffer[73]*(187))+$signed(in_buffer[74]*(188))+$signed(in_buffer[75]*(210));
assign in_buffer_weight42=$signed(in_buffer[50]*(41))+$signed(in_buffer[51]*(109))+$signed(in_buffer[52]*(108))+$signed(in_buffer[62]*(-58))+$signed(in_buffer[63]*(281))+$signed(in_buffer[64]*(143))+$signed(in_buffer[74]*(187))+$signed(in_buffer[75]*(188))+$signed(in_buffer[76]*(210));
assign in_buffer_weight43=$signed(in_buffer[51]*(41))+$signed(in_buffer[52]*(109))+$signed(in_buffer[53]*(108))+$signed(in_buffer[63]*(-58))+$signed(in_buffer[64]*(281))+$signed(in_buffer[65]*(143))+$signed(in_buffer[75]*(187))+$signed(in_buffer[76]*(188))+$signed(in_buffer[77]*(210));
assign in_buffer_weight44=$signed(in_buffer[52]*(41))+$signed(in_buffer[53]*(109))+$signed(in_buffer[54]*(108))+$signed(in_buffer[64]*(-58))+$signed(in_buffer[65]*(281))+$signed(in_buffer[66]*(143))+$signed(in_buffer[76]*(187))+$signed(in_buffer[77]*(188))+$signed(in_buffer[78]*(210));
assign in_buffer_weight45=$signed(in_buffer[53]*(41))+$signed(in_buffer[54]*(109))+$signed(in_buffer[55]*(108))+$signed(in_buffer[65]*(-58))+$signed(in_buffer[66]*(281))+$signed(in_buffer[67]*(143))+$signed(in_buffer[77]*(187))+$signed(in_buffer[78]*(188))+$signed(in_buffer[79]*(210));
assign in_buffer_weight46=$signed(in_buffer[54]*(41))+$signed(in_buffer[55]*(109))+$signed(in_buffer[56]*(108))+$signed(in_buffer[66]*(-58))+$signed(in_buffer[67]*(281))+$signed(in_buffer[68]*(143))+$signed(in_buffer[78]*(187))+$signed(in_buffer[79]*(188))+$signed(in_buffer[80]*(210));
assign in_buffer_weight47=$signed(in_buffer[55]*(41))+$signed(in_buffer[56]*(109))+$signed(in_buffer[57]*(108))+$signed(in_buffer[67]*(-58))+$signed(in_buffer[68]*(281))+$signed(in_buffer[69]*(143))+$signed(in_buffer[79]*(187))+$signed(in_buffer[80]*(188))+$signed(in_buffer[81]*(210));
assign in_buffer_weight48=$signed(in_buffer[56]*(41))+$signed(in_buffer[57]*(109))+$signed(in_buffer[58]*(108))+$signed(in_buffer[68]*(-58))+$signed(in_buffer[69]*(281))+$signed(in_buffer[70]*(143))+$signed(in_buffer[80]*(187))+$signed(in_buffer[81]*(188))+$signed(in_buffer[82]*(210));
assign in_buffer_weight49=$signed(in_buffer[57]*(41))+$signed(in_buffer[58]*(109))+$signed(in_buffer[59]*(108))+$signed(in_buffer[69]*(-58))+$signed(in_buffer[70]*(281))+$signed(in_buffer[71]*(143))+$signed(in_buffer[81]*(187))+$signed(in_buffer[82]*(188))+$signed(in_buffer[83]*(210));
assign in_buffer_weight50=$signed(in_buffer[60]*(41))+$signed(in_buffer[61]*(109))+$signed(in_buffer[62]*(108))+$signed(in_buffer[72]*(-58))+$signed(in_buffer[73]*(281))+$signed(in_buffer[74]*(143))+$signed(in_buffer[84]*(187))+$signed(in_buffer[85]*(188))+$signed(in_buffer[86]*(210));
assign in_buffer_weight51=$signed(in_buffer[61]*(41))+$signed(in_buffer[62]*(109))+$signed(in_buffer[63]*(108))+$signed(in_buffer[73]*(-58))+$signed(in_buffer[74]*(281))+$signed(in_buffer[75]*(143))+$signed(in_buffer[85]*(187))+$signed(in_buffer[86]*(188))+$signed(in_buffer[87]*(210));
assign in_buffer_weight52=$signed(in_buffer[62]*(41))+$signed(in_buffer[63]*(109))+$signed(in_buffer[64]*(108))+$signed(in_buffer[74]*(-58))+$signed(in_buffer[75]*(281))+$signed(in_buffer[76]*(143))+$signed(in_buffer[86]*(187))+$signed(in_buffer[87]*(188))+$signed(in_buffer[88]*(210));
assign in_buffer_weight53=$signed(in_buffer[63]*(41))+$signed(in_buffer[64]*(109))+$signed(in_buffer[65]*(108))+$signed(in_buffer[75]*(-58))+$signed(in_buffer[76]*(281))+$signed(in_buffer[77]*(143))+$signed(in_buffer[87]*(187))+$signed(in_buffer[88]*(188))+$signed(in_buffer[89]*(210));
assign in_buffer_weight54=$signed(in_buffer[64]*(41))+$signed(in_buffer[65]*(109))+$signed(in_buffer[66]*(108))+$signed(in_buffer[76]*(-58))+$signed(in_buffer[77]*(281))+$signed(in_buffer[78]*(143))+$signed(in_buffer[88]*(187))+$signed(in_buffer[89]*(188))+$signed(in_buffer[90]*(210));
assign in_buffer_weight55=$signed(in_buffer[65]*(41))+$signed(in_buffer[66]*(109))+$signed(in_buffer[67]*(108))+$signed(in_buffer[77]*(-58))+$signed(in_buffer[78]*(281))+$signed(in_buffer[79]*(143))+$signed(in_buffer[89]*(187))+$signed(in_buffer[90]*(188))+$signed(in_buffer[91]*(210));
assign in_buffer_weight56=$signed(in_buffer[66]*(41))+$signed(in_buffer[67]*(109))+$signed(in_buffer[68]*(108))+$signed(in_buffer[78]*(-58))+$signed(in_buffer[79]*(281))+$signed(in_buffer[80]*(143))+$signed(in_buffer[90]*(187))+$signed(in_buffer[91]*(188))+$signed(in_buffer[92]*(210));
assign in_buffer_weight57=$signed(in_buffer[67]*(41))+$signed(in_buffer[68]*(109))+$signed(in_buffer[69]*(108))+$signed(in_buffer[79]*(-58))+$signed(in_buffer[80]*(281))+$signed(in_buffer[81]*(143))+$signed(in_buffer[91]*(187))+$signed(in_buffer[92]*(188))+$signed(in_buffer[93]*(210));
assign in_buffer_weight58=$signed(in_buffer[68]*(41))+$signed(in_buffer[69]*(109))+$signed(in_buffer[70]*(108))+$signed(in_buffer[80]*(-58))+$signed(in_buffer[81]*(281))+$signed(in_buffer[82]*(143))+$signed(in_buffer[92]*(187))+$signed(in_buffer[93]*(188))+$signed(in_buffer[94]*(210));
assign in_buffer_weight59=$signed(in_buffer[69]*(41))+$signed(in_buffer[70]*(109))+$signed(in_buffer[71]*(108))+$signed(in_buffer[81]*(-58))+$signed(in_buffer[82]*(281))+$signed(in_buffer[83]*(143))+$signed(in_buffer[93]*(187))+$signed(in_buffer[94]*(188))+$signed(in_buffer[95]*(210));
assign in_buffer_weight60=$signed(in_buffer[72]*(41))+$signed(in_buffer[73]*(109))+$signed(in_buffer[74]*(108))+$signed(in_buffer[84]*(-58))+$signed(in_buffer[85]*(281))+$signed(in_buffer[86]*(143))+$signed(in_buffer[96]*(187))+$signed(in_buffer[97]*(188))+$signed(in_buffer[98]*(210));
assign in_buffer_weight61=$signed(in_buffer[73]*(41))+$signed(in_buffer[74]*(109))+$signed(in_buffer[75]*(108))+$signed(in_buffer[85]*(-58))+$signed(in_buffer[86]*(281))+$signed(in_buffer[87]*(143))+$signed(in_buffer[97]*(187))+$signed(in_buffer[98]*(188))+$signed(in_buffer[99]*(210));
assign in_buffer_weight62=$signed(in_buffer[74]*(41))+$signed(in_buffer[75]*(109))+$signed(in_buffer[76]*(108))+$signed(in_buffer[86]*(-58))+$signed(in_buffer[87]*(281))+$signed(in_buffer[88]*(143))+$signed(in_buffer[98]*(187))+$signed(in_buffer[99]*(188))+$signed(in_buffer[100]*(210));
assign in_buffer_weight63=$signed(in_buffer[75]*(41))+$signed(in_buffer[76]*(109))+$signed(in_buffer[77]*(108))+$signed(in_buffer[87]*(-58))+$signed(in_buffer[88]*(281))+$signed(in_buffer[89]*(143))+$signed(in_buffer[99]*(187))+$signed(in_buffer[100]*(188))+$signed(in_buffer[101]*(210));
assign in_buffer_weight64=$signed(in_buffer[76]*(41))+$signed(in_buffer[77]*(109))+$signed(in_buffer[78]*(108))+$signed(in_buffer[88]*(-58))+$signed(in_buffer[89]*(281))+$signed(in_buffer[90]*(143))+$signed(in_buffer[100]*(187))+$signed(in_buffer[101]*(188))+$signed(in_buffer[102]*(210));
assign in_buffer_weight65=$signed(in_buffer[77]*(41))+$signed(in_buffer[78]*(109))+$signed(in_buffer[79]*(108))+$signed(in_buffer[89]*(-58))+$signed(in_buffer[90]*(281))+$signed(in_buffer[91]*(143))+$signed(in_buffer[101]*(187))+$signed(in_buffer[102]*(188))+$signed(in_buffer[103]*(210));
assign in_buffer_weight66=$signed(in_buffer[78]*(41))+$signed(in_buffer[79]*(109))+$signed(in_buffer[80]*(108))+$signed(in_buffer[90]*(-58))+$signed(in_buffer[91]*(281))+$signed(in_buffer[92]*(143))+$signed(in_buffer[102]*(187))+$signed(in_buffer[103]*(188))+$signed(in_buffer[104]*(210));
assign in_buffer_weight67=$signed(in_buffer[79]*(41))+$signed(in_buffer[80]*(109))+$signed(in_buffer[81]*(108))+$signed(in_buffer[91]*(-58))+$signed(in_buffer[92]*(281))+$signed(in_buffer[93]*(143))+$signed(in_buffer[103]*(187))+$signed(in_buffer[104]*(188))+$signed(in_buffer[105]*(210));
assign in_buffer_weight68=$signed(in_buffer[80]*(41))+$signed(in_buffer[81]*(109))+$signed(in_buffer[82]*(108))+$signed(in_buffer[92]*(-58))+$signed(in_buffer[93]*(281))+$signed(in_buffer[94]*(143))+$signed(in_buffer[104]*(187))+$signed(in_buffer[105]*(188))+$signed(in_buffer[106]*(210));
assign in_buffer_weight69=$signed(in_buffer[81]*(41))+$signed(in_buffer[82]*(109))+$signed(in_buffer[83]*(108))+$signed(in_buffer[93]*(-58))+$signed(in_buffer[94]*(281))+$signed(in_buffer[95]*(143))+$signed(in_buffer[105]*(187))+$signed(in_buffer[106]*(188))+$signed(in_buffer[107]*(210));
assign in_buffer_weight70=$signed(in_buffer[84]*(41))+$signed(in_buffer[85]*(109))+$signed(in_buffer[86]*(108))+$signed(in_buffer[96]*(-58))+$signed(in_buffer[97]*(281))+$signed(in_buffer[98]*(143))+$signed(in_buffer[108]*(187))+$signed(in_buffer[109]*(188))+$signed(in_buffer[110]*(210));
assign in_buffer_weight71=$signed(in_buffer[85]*(41))+$signed(in_buffer[86]*(109))+$signed(in_buffer[87]*(108))+$signed(in_buffer[97]*(-58))+$signed(in_buffer[98]*(281))+$signed(in_buffer[99]*(143))+$signed(in_buffer[109]*(187))+$signed(in_buffer[110]*(188))+$signed(in_buffer[111]*(210));
assign in_buffer_weight72=$signed(in_buffer[86]*(41))+$signed(in_buffer[87]*(109))+$signed(in_buffer[88]*(108))+$signed(in_buffer[98]*(-58))+$signed(in_buffer[99]*(281))+$signed(in_buffer[100]*(143))+$signed(in_buffer[110]*(187))+$signed(in_buffer[111]*(188))+$signed(in_buffer[112]*(210));
assign in_buffer_weight73=$signed(in_buffer[87]*(41))+$signed(in_buffer[88]*(109))+$signed(in_buffer[89]*(108))+$signed(in_buffer[99]*(-58))+$signed(in_buffer[100]*(281))+$signed(in_buffer[101]*(143))+$signed(in_buffer[111]*(187))+$signed(in_buffer[112]*(188))+$signed(in_buffer[113]*(210));
assign in_buffer_weight74=$signed(in_buffer[88]*(41))+$signed(in_buffer[89]*(109))+$signed(in_buffer[90]*(108))+$signed(in_buffer[100]*(-58))+$signed(in_buffer[101]*(281))+$signed(in_buffer[102]*(143))+$signed(in_buffer[112]*(187))+$signed(in_buffer[113]*(188))+$signed(in_buffer[114]*(210));
assign in_buffer_weight75=$signed(in_buffer[89]*(41))+$signed(in_buffer[90]*(109))+$signed(in_buffer[91]*(108))+$signed(in_buffer[101]*(-58))+$signed(in_buffer[102]*(281))+$signed(in_buffer[103]*(143))+$signed(in_buffer[113]*(187))+$signed(in_buffer[114]*(188))+$signed(in_buffer[115]*(210));
assign in_buffer_weight76=$signed(in_buffer[90]*(41))+$signed(in_buffer[91]*(109))+$signed(in_buffer[92]*(108))+$signed(in_buffer[102]*(-58))+$signed(in_buffer[103]*(281))+$signed(in_buffer[104]*(143))+$signed(in_buffer[114]*(187))+$signed(in_buffer[115]*(188))+$signed(in_buffer[116]*(210));
assign in_buffer_weight77=$signed(in_buffer[91]*(41))+$signed(in_buffer[92]*(109))+$signed(in_buffer[93]*(108))+$signed(in_buffer[103]*(-58))+$signed(in_buffer[104]*(281))+$signed(in_buffer[105]*(143))+$signed(in_buffer[115]*(187))+$signed(in_buffer[116]*(188))+$signed(in_buffer[117]*(210));
assign in_buffer_weight78=$signed(in_buffer[92]*(41))+$signed(in_buffer[93]*(109))+$signed(in_buffer[94]*(108))+$signed(in_buffer[104]*(-58))+$signed(in_buffer[105]*(281))+$signed(in_buffer[106]*(143))+$signed(in_buffer[116]*(187))+$signed(in_buffer[117]*(188))+$signed(in_buffer[118]*(210));
assign in_buffer_weight79=$signed(in_buffer[93]*(41))+$signed(in_buffer[94]*(109))+$signed(in_buffer[95]*(108))+$signed(in_buffer[105]*(-58))+$signed(in_buffer[106]*(281))+$signed(in_buffer[107]*(143))+$signed(in_buffer[117]*(187))+$signed(in_buffer[118]*(188))+$signed(in_buffer[119]*(210));
assign in_buffer_weight80=$signed(in_buffer[96]*(41))+$signed(in_buffer[97]*(109))+$signed(in_buffer[98]*(108))+$signed(in_buffer[108]*(-58))+$signed(in_buffer[109]*(281))+$signed(in_buffer[110]*(143))+$signed(in_buffer[120]*(187))+$signed(in_buffer[121]*(188))+$signed(in_buffer[122]*(210));
assign in_buffer_weight81=$signed(in_buffer[97]*(41))+$signed(in_buffer[98]*(109))+$signed(in_buffer[99]*(108))+$signed(in_buffer[109]*(-58))+$signed(in_buffer[110]*(281))+$signed(in_buffer[111]*(143))+$signed(in_buffer[121]*(187))+$signed(in_buffer[122]*(188))+$signed(in_buffer[123]*(210));
assign in_buffer_weight82=$signed(in_buffer[98]*(41))+$signed(in_buffer[99]*(109))+$signed(in_buffer[100]*(108))+$signed(in_buffer[110]*(-58))+$signed(in_buffer[111]*(281))+$signed(in_buffer[112]*(143))+$signed(in_buffer[122]*(187))+$signed(in_buffer[123]*(188))+$signed(in_buffer[124]*(210));
assign in_buffer_weight83=$signed(in_buffer[99]*(41))+$signed(in_buffer[100]*(109))+$signed(in_buffer[101]*(108))+$signed(in_buffer[111]*(-58))+$signed(in_buffer[112]*(281))+$signed(in_buffer[113]*(143))+$signed(in_buffer[123]*(187))+$signed(in_buffer[124]*(188))+$signed(in_buffer[125]*(210));
assign in_buffer_weight84=$signed(in_buffer[100]*(41))+$signed(in_buffer[101]*(109))+$signed(in_buffer[102]*(108))+$signed(in_buffer[112]*(-58))+$signed(in_buffer[113]*(281))+$signed(in_buffer[114]*(143))+$signed(in_buffer[124]*(187))+$signed(in_buffer[125]*(188))+$signed(in_buffer[126]*(210));
assign in_buffer_weight85=$signed(in_buffer[101]*(41))+$signed(in_buffer[102]*(109))+$signed(in_buffer[103]*(108))+$signed(in_buffer[113]*(-58))+$signed(in_buffer[114]*(281))+$signed(in_buffer[115]*(143))+$signed(in_buffer[125]*(187))+$signed(in_buffer[126]*(188))+$signed(in_buffer[127]*(210));
assign in_buffer_weight86=$signed(in_buffer[102]*(41))+$signed(in_buffer[103]*(109))+$signed(in_buffer[104]*(108))+$signed(in_buffer[114]*(-58))+$signed(in_buffer[115]*(281))+$signed(in_buffer[116]*(143))+$signed(in_buffer[126]*(187))+$signed(in_buffer[127]*(188))+$signed(in_buffer[128]*(210));
assign in_buffer_weight87=$signed(in_buffer[103]*(41))+$signed(in_buffer[104]*(109))+$signed(in_buffer[105]*(108))+$signed(in_buffer[115]*(-58))+$signed(in_buffer[116]*(281))+$signed(in_buffer[117]*(143))+$signed(in_buffer[127]*(187))+$signed(in_buffer[128]*(188))+$signed(in_buffer[129]*(210));
assign in_buffer_weight88=$signed(in_buffer[104]*(41))+$signed(in_buffer[105]*(109))+$signed(in_buffer[106]*(108))+$signed(in_buffer[116]*(-58))+$signed(in_buffer[117]*(281))+$signed(in_buffer[118]*(143))+$signed(in_buffer[128]*(187))+$signed(in_buffer[129]*(188))+$signed(in_buffer[130]*(210));
assign in_buffer_weight89=$signed(in_buffer[105]*(41))+$signed(in_buffer[106]*(109))+$signed(in_buffer[107]*(108))+$signed(in_buffer[117]*(-58))+$signed(in_buffer[118]*(281))+$signed(in_buffer[119]*(143))+$signed(in_buffer[129]*(187))+$signed(in_buffer[130]*(188))+$signed(in_buffer[131]*(210));
assign in_buffer_weight90=$signed(in_buffer[108]*(41))+$signed(in_buffer[109]*(109))+$signed(in_buffer[110]*(108))+$signed(in_buffer[120]*(-58))+$signed(in_buffer[121]*(281))+$signed(in_buffer[122]*(143))+$signed(in_buffer[132]*(187))+$signed(in_buffer[133]*(188))+$signed(in_buffer[134]*(210));
assign in_buffer_weight91=$signed(in_buffer[109]*(41))+$signed(in_buffer[110]*(109))+$signed(in_buffer[111]*(108))+$signed(in_buffer[121]*(-58))+$signed(in_buffer[122]*(281))+$signed(in_buffer[123]*(143))+$signed(in_buffer[133]*(187))+$signed(in_buffer[134]*(188))+$signed(in_buffer[135]*(210));
assign in_buffer_weight92=$signed(in_buffer[110]*(41))+$signed(in_buffer[111]*(109))+$signed(in_buffer[112]*(108))+$signed(in_buffer[122]*(-58))+$signed(in_buffer[123]*(281))+$signed(in_buffer[124]*(143))+$signed(in_buffer[134]*(187))+$signed(in_buffer[135]*(188))+$signed(in_buffer[136]*(210));
assign in_buffer_weight93=$signed(in_buffer[111]*(41))+$signed(in_buffer[112]*(109))+$signed(in_buffer[113]*(108))+$signed(in_buffer[123]*(-58))+$signed(in_buffer[124]*(281))+$signed(in_buffer[125]*(143))+$signed(in_buffer[135]*(187))+$signed(in_buffer[136]*(188))+$signed(in_buffer[137]*(210));
assign in_buffer_weight94=$signed(in_buffer[112]*(41))+$signed(in_buffer[113]*(109))+$signed(in_buffer[114]*(108))+$signed(in_buffer[124]*(-58))+$signed(in_buffer[125]*(281))+$signed(in_buffer[126]*(143))+$signed(in_buffer[136]*(187))+$signed(in_buffer[137]*(188))+$signed(in_buffer[138]*(210));
assign in_buffer_weight95=$signed(in_buffer[113]*(41))+$signed(in_buffer[114]*(109))+$signed(in_buffer[115]*(108))+$signed(in_buffer[125]*(-58))+$signed(in_buffer[126]*(281))+$signed(in_buffer[127]*(143))+$signed(in_buffer[137]*(187))+$signed(in_buffer[138]*(188))+$signed(in_buffer[139]*(210));
assign in_buffer_weight96=$signed(in_buffer[114]*(41))+$signed(in_buffer[115]*(109))+$signed(in_buffer[116]*(108))+$signed(in_buffer[126]*(-58))+$signed(in_buffer[127]*(281))+$signed(in_buffer[128]*(143))+$signed(in_buffer[138]*(187))+$signed(in_buffer[139]*(188))+$signed(in_buffer[140]*(210));
assign in_buffer_weight97=$signed(in_buffer[115]*(41))+$signed(in_buffer[116]*(109))+$signed(in_buffer[117]*(108))+$signed(in_buffer[127]*(-58))+$signed(in_buffer[128]*(281))+$signed(in_buffer[129]*(143))+$signed(in_buffer[139]*(187))+$signed(in_buffer[140]*(188))+$signed(in_buffer[141]*(210));
assign in_buffer_weight98=$signed(in_buffer[116]*(41))+$signed(in_buffer[117]*(109))+$signed(in_buffer[118]*(108))+$signed(in_buffer[128]*(-58))+$signed(in_buffer[129]*(281))+$signed(in_buffer[130]*(143))+$signed(in_buffer[140]*(187))+$signed(in_buffer[141]*(188))+$signed(in_buffer[142]*(210));
assign in_buffer_weight99=$signed(in_buffer[117]*(41))+$signed(in_buffer[118]*(109))+$signed(in_buffer[119]*(108))+$signed(in_buffer[129]*(-58))+$signed(in_buffer[130]*(281))+$signed(in_buffer[131]*(143))+$signed(in_buffer[141]*(187))+$signed(in_buffer[142]*(188))+$signed(in_buffer[143]*(210));
wire signed    [DATA_WIDTH-1:0]   weight_bias0;
assign weight_bias0= in_buffer_weight0+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias1;
assign weight_bias1= in_buffer_weight1+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias2;
assign weight_bias2= in_buffer_weight2+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias3;
assign weight_bias3= in_buffer_weight3+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias4;
assign weight_bias4= in_buffer_weight4+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias5;
assign weight_bias5= in_buffer_weight5+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias6;
assign weight_bias6= in_buffer_weight6+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias7;
assign weight_bias7= in_buffer_weight7+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias8;
assign weight_bias8= in_buffer_weight8+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias9= in_buffer_weight9+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias10;
assign weight_bias10= in_buffer_weight10+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias11;
assign weight_bias11= in_buffer_weight11+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias12;
assign weight_bias12= in_buffer_weight12+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias13;
assign weight_bias13= in_buffer_weight13+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias14;
assign weight_bias14= in_buffer_weight14+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias15;
assign weight_bias15= in_buffer_weight15+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias16;
assign weight_bias16= in_buffer_weight16+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias17;
assign weight_bias17= in_buffer_weight17+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias18;
assign weight_bias18= in_buffer_weight18+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias19;
assign weight_bias19= in_buffer_weight19+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias20;
assign weight_bias20= in_buffer_weight20+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias21;
assign weight_bias21= in_buffer_weight21+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias22;
assign weight_bias22= in_buffer_weight22+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias23;
assign weight_bias23= in_buffer_weight23+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias24;
assign weight_bias24= in_buffer_weight24+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias25;
assign weight_bias25= in_buffer_weight25+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias26;
assign weight_bias26= in_buffer_weight26+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias27;
assign weight_bias27= in_buffer_weight27+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias28;
assign weight_bias28= in_buffer_weight28+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias29;
assign weight_bias29= in_buffer_weight29+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias30;
assign weight_bias30= in_buffer_weight30+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias31;
assign weight_bias31= in_buffer_weight31+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias32;
assign weight_bias32= in_buffer_weight32+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias33;
assign weight_bias33= in_buffer_weight33+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias34;
assign weight_bias34= in_buffer_weight34+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias35;
assign weight_bias35= in_buffer_weight35+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias36;
assign weight_bias36= in_buffer_weight36+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias37;
assign weight_bias37= in_buffer_weight37+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias38;
assign weight_bias38= in_buffer_weight38+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias39;
assign weight_bias39= in_buffer_weight39+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias40;
assign weight_bias40= in_buffer_weight40+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias41;
assign weight_bias41= in_buffer_weight41+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias42;
assign weight_bias42= in_buffer_weight42+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias43;
assign weight_bias43= in_buffer_weight43+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias44;
assign weight_bias44= in_buffer_weight44+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias45;
assign weight_bias45= in_buffer_weight45+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias46;
assign weight_bias46= in_buffer_weight46+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias47;
assign weight_bias47= in_buffer_weight47+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias48;
assign weight_bias48= in_buffer_weight48+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias49;
assign weight_bias49= in_buffer_weight49+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias50;
assign weight_bias50= in_buffer_weight50+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias51;
assign weight_bias51= in_buffer_weight51+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias52;
assign weight_bias52= in_buffer_weight52+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias53;
assign weight_bias53= in_buffer_weight53+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias54;
assign weight_bias54= in_buffer_weight54+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias55;
assign weight_bias55= in_buffer_weight55+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias56;
assign weight_bias56= in_buffer_weight56+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias57;
assign weight_bias57= in_buffer_weight57+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias58;
assign weight_bias58= in_buffer_weight58+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias59;
assign weight_bias59= in_buffer_weight59+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias60;
assign weight_bias60= in_buffer_weight60+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias61;
assign weight_bias61= in_buffer_weight61+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias62;
assign weight_bias62= in_buffer_weight62+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias63;
assign weight_bias63= in_buffer_weight63+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias64;
assign weight_bias64= in_buffer_weight64+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias65;
assign weight_bias65= in_buffer_weight65+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias66;
assign weight_bias66= in_buffer_weight66+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias67;
assign weight_bias67= in_buffer_weight67+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias68;
assign weight_bias68= in_buffer_weight68+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias69;
assign weight_bias69= in_buffer_weight69+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias70;
assign weight_bias70= in_buffer_weight70+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias71;
assign weight_bias71= in_buffer_weight71+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias72;
assign weight_bias72= in_buffer_weight72+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias73;
assign weight_bias73= in_buffer_weight73+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias74;
assign weight_bias74= in_buffer_weight74+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias75;
assign weight_bias75= in_buffer_weight75+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias76;
assign weight_bias76= in_buffer_weight76+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias77;
assign weight_bias77= in_buffer_weight77+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias78;
assign weight_bias78= in_buffer_weight78+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias79;
assign weight_bias79= in_buffer_weight79+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias80;
assign weight_bias80= in_buffer_weight80+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias81;
assign weight_bias81= in_buffer_weight81+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias82;
assign weight_bias82= in_buffer_weight82+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias83;
assign weight_bias83= in_buffer_weight83+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias84;
assign weight_bias84= in_buffer_weight84+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias85;
assign weight_bias85= in_buffer_weight85+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias86;
assign weight_bias86= in_buffer_weight86+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias87;
assign weight_bias87= in_buffer_weight87+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias88;
assign weight_bias88= in_buffer_weight88+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias89;
assign weight_bias89= in_buffer_weight89+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias90;
assign weight_bias90= in_buffer_weight90+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias91;
assign weight_bias91= in_buffer_weight91+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias92;
assign weight_bias92= in_buffer_weight92+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias93;
assign weight_bias93= in_buffer_weight93+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias94;
assign weight_bias94= in_buffer_weight94+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias95;
assign weight_bias95= in_buffer_weight95+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias96;
assign weight_bias96= in_buffer_weight96+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias97;
assign weight_bias97= in_buffer_weight97+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias98;
assign weight_bias98= in_buffer_weight98+0;
wire signed    [DATA_WIDTH-1:0]   weight_bias99;
assign weight_bias99= in_buffer_weight99+0;
wire signed    [DATA_WIDTH-1:0]   bias_relu0;
wire signed    [DATA_WIDTH-1:0]   bias_relu1;
wire signed    [DATA_WIDTH-1:0]   bias_relu2;
wire signed    [DATA_WIDTH-1:0]   bias_relu3;
wire signed    [DATA_WIDTH-1:0]   bias_relu4;
wire signed    [DATA_WIDTH-1:0]   bias_relu5;
wire signed    [DATA_WIDTH-1:0]   bias_relu6;
wire signed    [DATA_WIDTH-1:0]   bias_relu7;
wire signed    [DATA_WIDTH-1:0]   bias_relu8;
wire signed    [DATA_WIDTH-1:0]   bias_relu9;
wire signed    [DATA_WIDTH-1:0]   bias_relu10;
wire signed    [DATA_WIDTH-1:0]   bias_relu11;
wire signed    [DATA_WIDTH-1:0]   bias_relu12;
wire signed    [DATA_WIDTH-1:0]   bias_relu13;
wire signed    [DATA_WIDTH-1:0]   bias_relu14;
wire signed    [DATA_WIDTH-1:0]   bias_relu15;
wire signed    [DATA_WIDTH-1:0]   bias_relu16;
wire signed    [DATA_WIDTH-1:0]   bias_relu17;
wire signed    [DATA_WIDTH-1:0]   bias_relu18;
wire signed    [DATA_WIDTH-1:0]   bias_relu19;
wire signed    [DATA_WIDTH-1:0]   bias_relu20;
wire signed    [DATA_WIDTH-1:0]   bias_relu21;
wire signed    [DATA_WIDTH-1:0]   bias_relu22;
wire signed    [DATA_WIDTH-1:0]   bias_relu23;
wire signed    [DATA_WIDTH-1:0]   bias_relu24;
wire signed    [DATA_WIDTH-1:0]   bias_relu25;
wire signed    [DATA_WIDTH-1:0]   bias_relu26;
wire signed    [DATA_WIDTH-1:0]   bias_relu27;
wire signed    [DATA_WIDTH-1:0]   bias_relu28;
wire signed    [DATA_WIDTH-1:0]   bias_relu29;
wire signed    [DATA_WIDTH-1:0]   bias_relu30;
wire signed    [DATA_WIDTH-1:0]   bias_relu31;
wire signed    [DATA_WIDTH-1:0]   bias_relu32;
wire signed    [DATA_WIDTH-1:0]   bias_relu33;
wire signed    [DATA_WIDTH-1:0]   bias_relu34;
wire signed    [DATA_WIDTH-1:0]   bias_relu35;
wire signed    [DATA_WIDTH-1:0]   bias_relu36;
wire signed    [DATA_WIDTH-1:0]   bias_relu37;
wire signed    [DATA_WIDTH-1:0]   bias_relu38;
wire signed    [DATA_WIDTH-1:0]   bias_relu39;
wire signed    [DATA_WIDTH-1:0]   bias_relu40;
wire signed    [DATA_WIDTH-1:0]   bias_relu41;
wire signed    [DATA_WIDTH-1:0]   bias_relu42;
wire signed    [DATA_WIDTH-1:0]   bias_relu43;
wire signed    [DATA_WIDTH-1:0]   bias_relu44;
wire signed    [DATA_WIDTH-1:0]   bias_relu45;
wire signed    [DATA_WIDTH-1:0]   bias_relu46;
wire signed    [DATA_WIDTH-1:0]   bias_relu47;
wire signed    [DATA_WIDTH-1:0]   bias_relu48;
wire signed    [DATA_WIDTH-1:0]   bias_relu49;
wire signed    [DATA_WIDTH-1:0]   bias_relu50;
wire signed    [DATA_WIDTH-1:0]   bias_relu51;
wire signed    [DATA_WIDTH-1:0]   bias_relu52;
wire signed    [DATA_WIDTH-1:0]   bias_relu53;
wire signed    [DATA_WIDTH-1:0]   bias_relu54;
wire signed    [DATA_WIDTH-1:0]   bias_relu55;
wire signed    [DATA_WIDTH-1:0]   bias_relu56;
wire signed    [DATA_WIDTH-1:0]   bias_relu57;
wire signed    [DATA_WIDTH-1:0]   bias_relu58;
wire signed    [DATA_WIDTH-1:0]   bias_relu59;
wire signed    [DATA_WIDTH-1:0]   bias_relu60;
wire signed    [DATA_WIDTH-1:0]   bias_relu61;
wire signed    [DATA_WIDTH-1:0]   bias_relu62;
wire signed    [DATA_WIDTH-1:0]   bias_relu63;
wire signed    [DATA_WIDTH-1:0]   bias_relu64;
wire signed    [DATA_WIDTH-1:0]   bias_relu65;
wire signed    [DATA_WIDTH-1:0]   bias_relu66;
wire signed    [DATA_WIDTH-1:0]   bias_relu67;
wire signed    [DATA_WIDTH-1:0]   bias_relu68;
wire signed    [DATA_WIDTH-1:0]   bias_relu69;
wire signed    [DATA_WIDTH-1:0]   bias_relu70;
wire signed    [DATA_WIDTH-1:0]   bias_relu71;
wire signed    [DATA_WIDTH-1:0]   bias_relu72;
wire signed    [DATA_WIDTH-1:0]   bias_relu73;
wire signed    [DATA_WIDTH-1:0]   bias_relu74;
wire signed    [DATA_WIDTH-1:0]   bias_relu75;
wire signed    [DATA_WIDTH-1:0]   bias_relu76;
wire signed    [DATA_WIDTH-1:0]   bias_relu77;
wire signed    [DATA_WIDTH-1:0]   bias_relu78;
wire signed    [DATA_WIDTH-1:0]   bias_relu79;
wire signed    [DATA_WIDTH-1:0]   bias_relu80;
wire signed    [DATA_WIDTH-1:0]   bias_relu81;
wire signed    [DATA_WIDTH-1:0]   bias_relu82;
wire signed    [DATA_WIDTH-1:0]   bias_relu83;
wire signed    [DATA_WIDTH-1:0]   bias_relu84;
wire signed    [DATA_WIDTH-1:0]   bias_relu85;
wire signed    [DATA_WIDTH-1:0]   bias_relu86;
wire signed    [DATA_WIDTH-1:0]   bias_relu87;
wire signed    [DATA_WIDTH-1:0]   bias_relu88;
wire signed    [DATA_WIDTH-1:0]   bias_relu89;
wire signed    [DATA_WIDTH-1:0]   bias_relu90;
wire signed    [DATA_WIDTH-1:0]   bias_relu91;
wire signed    [DATA_WIDTH-1:0]   bias_relu92;
wire signed    [DATA_WIDTH-1:0]   bias_relu93;
wire signed    [DATA_WIDTH-1:0]   bias_relu94;
wire signed    [DATA_WIDTH-1:0]   bias_relu95;
wire signed    [DATA_WIDTH-1:0]   bias_relu96;
wire signed    [DATA_WIDTH-1:0]   bias_relu97;
wire signed    [DATA_WIDTH-1:0]   bias_relu98;
wire signed    [DATA_WIDTH-1:0]   bias_relu99;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign bias_relu32=(weight_bias32[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias32;
assign bias_relu33=(weight_bias33[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias33;
assign bias_relu34=(weight_bias34[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias34;
assign bias_relu35=(weight_bias35[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias35;
assign bias_relu36=(weight_bias36[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias36;
assign bias_relu37=(weight_bias37[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias37;
assign bias_relu38=(weight_bias38[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias38;
assign bias_relu39=(weight_bias39[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias39;
assign bias_relu40=(weight_bias40[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias40;
assign bias_relu41=(weight_bias41[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias41;
assign bias_relu42=(weight_bias42[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias42;
assign bias_relu43=(weight_bias43[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias43;
assign bias_relu44=(weight_bias44[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias44;
assign bias_relu45=(weight_bias45[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias45;
assign bias_relu46=(weight_bias46[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias46;
assign bias_relu47=(weight_bias47[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias47;
assign bias_relu48=(weight_bias48[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias48;
assign bias_relu49=(weight_bias49[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias49;
assign bias_relu50=(weight_bias50[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias50;
assign bias_relu51=(weight_bias51[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias51;
assign bias_relu52=(weight_bias52[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias52;
assign bias_relu53=(weight_bias53[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias53;
assign bias_relu54=(weight_bias54[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias54;
assign bias_relu55=(weight_bias55[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias55;
assign bias_relu56=(weight_bias56[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias56;
assign bias_relu57=(weight_bias57[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias57;
assign bias_relu58=(weight_bias58[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias58;
assign bias_relu59=(weight_bias59[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias59;
assign bias_relu60=(weight_bias60[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias60;
assign bias_relu61=(weight_bias61[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias61;
assign bias_relu62=(weight_bias62[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias62;
assign bias_relu63=(weight_bias63[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias63;
assign bias_relu64=(weight_bias64[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias64;
assign bias_relu65=(weight_bias65[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias65;
assign bias_relu66=(weight_bias66[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias66;
assign bias_relu67=(weight_bias67[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias67;
assign bias_relu68=(weight_bias68[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias68;
assign bias_relu69=(weight_bias69[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias69;
assign bias_relu70=(weight_bias70[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias70;
assign bias_relu71=(weight_bias71[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias71;
assign bias_relu72=(weight_bias72[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias72;
assign bias_relu73=(weight_bias73[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias73;
assign bias_relu74=(weight_bias74[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias74;
assign bias_relu75=(weight_bias75[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias75;
assign bias_relu76=(weight_bias76[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias76;
assign bias_relu77=(weight_bias77[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias77;
assign bias_relu78=(weight_bias78[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias78;
assign bias_relu79=(weight_bias79[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias79;
assign bias_relu80=(weight_bias80[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias80;
assign bias_relu81=(weight_bias81[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias81;
assign bias_relu82=(weight_bias82[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias82;
assign bias_relu83=(weight_bias83[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias83;
assign bias_relu84=(weight_bias84[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias84;
assign bias_relu85=(weight_bias85[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias85;
assign bias_relu86=(weight_bias86[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias86;
assign bias_relu87=(weight_bias87[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias87;
assign bias_relu88=(weight_bias88[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias88;
assign bias_relu89=(weight_bias89[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias89;
assign bias_relu90=(weight_bias90[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias90;
assign bias_relu91=(weight_bias91[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias91;
assign bias_relu92=(weight_bias92[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias92;
assign bias_relu93=(weight_bias93[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias93;
assign bias_relu94=(weight_bias94[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias94;
assign bias_relu95=(weight_bias95[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias95;
assign bias_relu96=(weight_bias96[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias96;
assign bias_relu97=(weight_bias97[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias97;
assign bias_relu98=(weight_bias98[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias98;
assign bias_relu99=(weight_bias99[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias99;
always@(posedge clk)
    begin
        if(~rst)
            begin
           layer_out <={bias_relu99,bias_relu98,bias_relu97,bias_relu96,bias_relu95,bias_relu94,bias_relu93,bias_relu92,bias_relu91,bias_relu90,bias_relu89,bias_relu88,bias_relu87,bias_relu86,bias_relu85,bias_relu84,bias_relu83,bias_relu82,bias_relu81,bias_relu80,bias_relu79,bias_relu78,bias_relu77,bias_relu76,bias_relu75,bias_relu74,bias_relu73,bias_relu72,bias_relu71,bias_relu70,bias_relu69,bias_relu68,bias_relu67,bias_relu66,bias_relu65,bias_relu64,bias_relu63,bias_relu62,bias_relu61,bias_relu60,bias_relu59,bias_relu58,bias_relu57,bias_relu56,bias_relu55,bias_relu54,bias_relu53,bias_relu52,bias_relu51,bias_relu50,bias_relu49,bias_relu48,bias_relu47,bias_relu46,bias_relu45,bias_relu44,bias_relu43,bias_relu42,bias_relu41,bias_relu40,bias_relu39,bias_relu38,bias_relu37,bias_relu36,bias_relu35,bias_relu34,bias_relu33,bias_relu32,bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
            end
        else
            begin
           layer_out<= {(OUTPUT_BIT*OUTPUT_NODE){1'b0}};
        end
    end
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule