module layer0_tcb_144x64x10
(
    input clk,
    input rst,
    input [144*8-1:0] img,
    input valid,
    output  reg ready,
    output [20*64-1:0] layer_out
);
parameter DATA_WIDTH = 20;
parameter IMG_SZ   =   144;
reg    signed [8-1:0]  in_buffer[0:IMG_SZ-1];
integer i;
always@(posedge clk )
    begin
        if(rst)
            begin
                for(i=0;i<IMG_SZ;i=i+1)
                    begin
                        in_buffer[i]<=0;
                    end
            end
        else
        begin
       in_buffer[0]<=img[7:0];
       in_buffer[1]<=img[15:8];
       in_buffer[2]<=img[23:16];
       in_buffer[3]<=img[31:24];
       in_buffer[4]<=img[39:32];
       in_buffer[5]<=img[47:40];
       in_buffer[6]<=img[55:48];
       in_buffer[7]<=img[63:56];
       in_buffer[8]<=img[71:64];
       in_buffer[9]<=img[79:72];
       in_buffer[10]<=img[87:80];
       in_buffer[11]<=img[95:88];
       in_buffer[12]<=img[103:96];
       in_buffer[13]<=img[111:104];
       in_buffer[14]<=img[119:112];
       in_buffer[15]<=img[127:120];
       in_buffer[16]<=img[135:128];
       in_buffer[17]<=img[143:136];
       in_buffer[18]<=img[151:144];
       in_buffer[19]<=img[159:152];
       in_buffer[20]<=img[167:160];
       in_buffer[21]<=img[175:168];
       in_buffer[22]<=img[183:176];
       in_buffer[23]<=img[191:184];
       in_buffer[24]<=img[199:192];
       in_buffer[25]<=img[207:200];
       in_buffer[26]<=img[215:208];
       in_buffer[27]<=img[223:216];
       in_buffer[28]<=img[231:224];
       in_buffer[29]<=img[239:232];
       in_buffer[30]<=img[247:240];
       in_buffer[31]<=img[255:248];
       in_buffer[32]<=img[263:256];
       in_buffer[33]<=img[271:264];
       in_buffer[34]<=img[279:272];
       in_buffer[35]<=img[287:280];
       in_buffer[36]<=img[295:288];
       in_buffer[37]<=img[303:296];
       in_buffer[38]<=img[311:304];
       in_buffer[39]<=img[319:312];
       in_buffer[40]<=img[327:320];
       in_buffer[41]<=img[335:328];
       in_buffer[42]<=img[343:336];
       in_buffer[43]<=img[351:344];
       in_buffer[44]<=img[359:352];
       in_buffer[45]<=img[367:360];
       in_buffer[46]<=img[375:368];
       in_buffer[47]<=img[383:376];
       in_buffer[48]<=img[391:384];
       in_buffer[49]<=img[399:392];
       in_buffer[50]<=img[407:400];
       in_buffer[51]<=img[415:408];
       in_buffer[52]<=img[423:416];
       in_buffer[53]<=img[431:424];
       in_buffer[54]<=img[439:432];
       in_buffer[55]<=img[447:440];
       in_buffer[56]<=img[455:448];
       in_buffer[57]<=img[463:456];
       in_buffer[58]<=img[471:464];
       in_buffer[59]<=img[479:472];
       in_buffer[60]<=img[487:480];
       in_buffer[61]<=img[495:488];
       in_buffer[62]<=img[503:496];
       in_buffer[63]<=img[511:504];
       in_buffer[64]<=img[519:512];
       in_buffer[65]<=img[527:520];
       in_buffer[66]<=img[535:528];
       in_buffer[67]<=img[543:536];
       in_buffer[68]<=img[551:544];
       in_buffer[69]<=img[559:552];
       in_buffer[70]<=img[567:560];
       in_buffer[71]<=img[575:568];
       in_buffer[72]<=img[583:576];
       in_buffer[73]<=img[591:584];
       in_buffer[74]<=img[599:592];
       in_buffer[75]<=img[607:600];
       in_buffer[76]<=img[615:608];
       in_buffer[77]<=img[623:616];
       in_buffer[78]<=img[631:624];
       in_buffer[79]<=img[639:632];
       in_buffer[80]<=img[647:640];
       in_buffer[81]<=img[655:648];
       in_buffer[82]<=img[663:656];
       in_buffer[83]<=img[671:664];
       in_buffer[84]<=img[679:672];
       in_buffer[85]<=img[687:680];
       in_buffer[86]<=img[695:688];
       in_buffer[87]<=img[703:696];
       in_buffer[88]<=img[711:704];
       in_buffer[89]<=img[719:712];
       in_buffer[90]<=img[727:720];
       in_buffer[91]<=img[735:728];
       in_buffer[92]<=img[743:736];
       in_buffer[93]<=img[751:744];
       in_buffer[94]<=img[759:752];
       in_buffer[95]<=img[767:760];
       in_buffer[96]<=img[775:768];
       in_buffer[97]<=img[783:776];
       in_buffer[98]<=img[791:784];
       in_buffer[99]<=img[799:792];
       in_buffer[100]<=img[807:800];
       in_buffer[101]<=img[815:808];
       in_buffer[102]<=img[823:816];
       in_buffer[103]<=img[831:824];
       in_buffer[104]<=img[839:832];
       in_buffer[105]<=img[847:840];
       in_buffer[106]<=img[855:848];
       in_buffer[107]<=img[863:856];
       in_buffer[108]<=img[871:864];
       in_buffer[109]<=img[879:872];
       in_buffer[110]<=img[887:880];
       in_buffer[111]<=img[895:888];
       in_buffer[112]<=img[903:896];
       in_buffer[113]<=img[911:904];
       in_buffer[114]<=img[919:912];
       in_buffer[115]<=img[927:920];
       in_buffer[116]<=img[935:928];
       in_buffer[117]<=img[943:936];
       in_buffer[118]<=img[951:944];
       in_buffer[119]<=img[959:952];
       in_buffer[120]<=img[967:960];
       in_buffer[121]<=img[975:968];
       in_buffer[122]<=img[983:976];
       in_buffer[123]<=img[991:984];
       in_buffer[124]<=img[999:992];
       in_buffer[125]<=img[1007:1000];
       in_buffer[126]<=img[1015:1008];
       in_buffer[127]<=img[1023:1016];
       in_buffer[128]<=img[1031:1024];
       in_buffer[129]<=img[1039:1032];
       in_buffer[130]<=img[1047:1040];
       in_buffer[131]<=img[1055:1048];
       in_buffer[132]<=img[1063:1056];
       in_buffer[133]<=img[1071:1064];
       in_buffer[134]<=img[1079:1072];
       in_buffer[135]<=img[1087:1080];
       in_buffer[136]<=img[1095:1088];
       in_buffer[137]<=img[1103:1096];
       in_buffer[138]<=img[1111:1104];
       in_buffer[139]<=img[1119:1112];
       in_buffer[140]<=img[1127:1120];
       in_buffer[141]<=img[1135:1128];
       in_buffer[142]<=img[1143:1136];
       in_buffer[143]<=img[1151:1144];
        end
   end
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0+(0-(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<6))+(0-(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<6))+(0-(in_buffer[9]<<0)-(in_buffer[9]<<2)+(in_buffer[9]<<6))+(0-(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<6))+(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<6))+(0-(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<6))+(0-(in_buffer[25]<<0)-(in_buffer[25]<<2)+(in_buffer[25]<<6))+(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)+(in_buffer[38]<<6))-(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))-(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))+(0-(in_buffer[46]<<0)-(in_buffer[46]<<2)+(in_buffer[46]<<6))+(0-(in_buffer[48]<<0)-(in_buffer[48]<<2)+(in_buffer[48]<<6))-(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<6))-(0-(in_buffer[109]<<0)-(in_buffer[109]<<2)+(in_buffer[109]<<6))-(0-(in_buffer[121]<<0)-(in_buffer[121]<<2)+(in_buffer[121]<<6))-(0-(in_buffer[130]<<0)-(in_buffer[130]<<2)+(in_buffer[130]<<6))-(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))-(0-(in_buffer[133]<<0)-(in_buffer[133]<<2)+(in_buffer[133]<<6))-(0-(in_buffer[134]<<0)-(in_buffer[134]<<2)+(in_buffer[134]<<6))-(0-(in_buffer[136]<<0)-(in_buffer[136]<<2)+(in_buffer[136]<<6))-(0-(in_buffer[137]<<0)-(in_buffer[137]<<2)+(in_buffer[137]<<6))-(0-(in_buffer[138]<<0)-(in_buffer[138]<<2)+(in_buffer[138]<<6))-(0-(in_buffer[139]<<0)-(in_buffer[139]<<2)+(in_buffer[139]<<6))-(0-(in_buffer[140]<<0)-(in_buffer[140]<<2)+(in_buffer[140]<<6))-(0-(in_buffer[141]<<0)-(in_buffer[141]<<2)+(in_buffer[141]<<6))-(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0-(0-(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<6))-(0-(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<6))+(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<6))+(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))-(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)+(in_buffer[36]<<6))-(0-(in_buffer[37]<<0)-(in_buffer[37]<<2)+(in_buffer[37]<<6))+(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))+(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)+(in_buffer[40]<<6))+(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))+(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))-(0-(in_buffer[46]<<0)-(in_buffer[46]<<2)+(in_buffer[46]<<6))-(0-(in_buffer[47]<<0)-(in_buffer[47]<<2)+(in_buffer[47]<<6))+(0-(in_buffer[61]<<0)-(in_buffer[61]<<2)+(in_buffer[61]<<6))+(0-(in_buffer[73]<<0)-(in_buffer[73]<<2)+(in_buffer[73]<<6))-(0-(in_buffer[88]<<0)-(in_buffer[88]<<2)+(in_buffer[88]<<6))-(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)+(in_buffer[90]<<6))-(0-(in_buffer[91]<<0)-(in_buffer[91]<<2)+(in_buffer[91]<<6))-(0-(in_buffer[105]<<0)-(in_buffer[105]<<2)+(in_buffer[105]<<6))+(0-(in_buffer[109]<<0)-(in_buffer[109]<<2)+(in_buffer[109]<<6))+(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<6))+(0-(in_buffer[121]<<0)-(in_buffer[121]<<2)+(in_buffer[121]<<6))+(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))+(0-(in_buffer[133]<<0)-(in_buffer[133]<<2)+(in_buffer[133]<<6))+(0-(in_buffer[135]<<0)-(in_buffer[135]<<2)+(in_buffer[135]<<6))+(0-(in_buffer[136]<<0)-(in_buffer[136]<<2)+(in_buffer[136]<<6))+(0-(in_buffer[137]<<0)-(in_buffer[137]<<2)+(in_buffer[137]<<6))+(0-(in_buffer[138]<<0)-(in_buffer[138]<<2)+(in_buffer[138]<<6))+(0-(in_buffer[139]<<0)-(in_buffer[139]<<2)+(in_buffer[139]<<6))+(0-(in_buffer[140]<<0)-(in_buffer[140]<<2)+(in_buffer[140]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0-(0-(in_buffer[4]<<0)-(in_buffer[4]<<2)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<6))-(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)+(in_buffer[7]<<6))-(0-(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<6))-(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<6))-(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)+(in_buffer[36]<<6))-(0-(in_buffer[37]<<0)-(in_buffer[37]<<2)+(in_buffer[37]<<6))-(0-(in_buffer[46]<<0)-(in_buffer[46]<<2)+(in_buffer[46]<<6))-(0-(in_buffer[48]<<0)-(in_buffer[48]<<2)+(in_buffer[48]<<6))-(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)+(in_buffer[49]<<6))-(0-(in_buffer[57]<<0)-(in_buffer[57]<<2)+(in_buffer[57]<<6))-(0-(in_buffer[58]<<0)-(in_buffer[58]<<2)+(in_buffer[58]<<6))-(0-(in_buffer[62]<<0)-(in_buffer[62]<<2)+(in_buffer[62]<<6))-(0-(in_buffer[63]<<0)-(in_buffer[63]<<2)+(in_buffer[63]<<6))-(0-(in_buffer[69]<<0)-(in_buffer[69]<<2)+(in_buffer[69]<<6))-(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)+(in_buffer[70]<<6))-(0-(in_buffer[72]<<0)-(in_buffer[72]<<2)+(in_buffer[72]<<6))-(0-(in_buffer[95]<<0)-(in_buffer[95]<<2)+(in_buffer[95]<<6))-(0-(in_buffer[126]<<0)-(in_buffer[126]<<2)+(in_buffer[126]<<6))-(0-(in_buffer[128]<<0)-(in_buffer[128]<<2)+(in_buffer[128]<<6))+(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight10;
assign in_buffer_weight10=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight11;
assign in_buffer_weight11=0-(0-(in_buffer[0]<<0)-(in_buffer[0]<<2)+(in_buffer[0]<<6))-(0-(in_buffer[1]<<0)-(in_buffer[1]<<2)+(in_buffer[1]<<6))-(0-(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<6))+(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<6))-(0-(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<6))+(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))+(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))+(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))+(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))+(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))+(0-(in_buffer[67]<<0)-(in_buffer[67]<<2)+(in_buffer[67]<<6))-(0-(in_buffer[73]<<0)-(in_buffer[73]<<2)+(in_buffer[73]<<6))+(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)+(in_buffer[75]<<6))+(0-(in_buffer[76]<<0)-(in_buffer[76]<<2)+(in_buffer[76]<<6))+(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<2)+(in_buffer[80]<<6))+(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)+(in_buffer[81]<<6))+(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6))-(0-(in_buffer[98]<<0)-(in_buffer[98]<<2)+(in_buffer[98]<<6))+(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))+(0-(in_buffer[134]<<0)-(in_buffer[134]<<2)+(in_buffer[134]<<6))+(0-(in_buffer[141]<<0)-(in_buffer[141]<<2)+(in_buffer[141]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight12;
assign in_buffer_weight12=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight13;
assign in_buffer_weight13=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight14;
assign in_buffer_weight14=0+(0-(in_buffer[26]<<0)-(in_buffer[26]<<2)+(in_buffer[26]<<6))+(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))+(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))+(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))-(0-(in_buffer[62]<<0)-(in_buffer[62]<<2)+(in_buffer[62]<<6))+(0-(in_buffer[76]<<0)-(in_buffer[76]<<2)+(in_buffer[76]<<6))+(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)+(in_buffer[77]<<6))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6))+(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))+(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)+(in_buffer[81]<<6))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<6))+(0-(in_buffer[87]<<0)-(in_buffer[87]<<2)+(in_buffer[87]<<6))+(0-(in_buffer[94]<<0)-(in_buffer[94]<<2)+(in_buffer[94]<<6))+(0-(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<6))-(0-(in_buffer[102]<<0)-(in_buffer[102]<<2)+(in_buffer[102]<<6))-(0-(in_buffer[103]<<0)-(in_buffer[103]<<2)+(in_buffer[103]<<6))+(0-(in_buffer[109]<<0)-(in_buffer[109]<<2)+(in_buffer[109]<<6))+(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<6))+(0-(in_buffer[121]<<0)-(in_buffer[121]<<2)+(in_buffer[121]<<6))-(0-(in_buffer[127]<<0)-(in_buffer[127]<<2)+(in_buffer[127]<<6))-(0-(in_buffer[134]<<0)-(in_buffer[134]<<2)+(in_buffer[134]<<6))-(0-(in_buffer[135]<<0)-(in_buffer[135]<<2)+(in_buffer[135]<<6))-(0-(in_buffer[140]<<0)-(in_buffer[140]<<2)+(in_buffer[140]<<6))-(0-(in_buffer[141]<<0)-(in_buffer[141]<<2)+(in_buffer[141]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight15;
assign in_buffer_weight15=0+(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)+(in_buffer[17]<<6))-(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))-(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))-(0-(in_buffer[67]<<0)-(in_buffer[67]<<2)+(in_buffer[67]<<6))+(0-(in_buffer[88]<<0)-(in_buffer[88]<<2)+(in_buffer[88]<<6))+(0-(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<6))-(0-(in_buffer[95]<<0)-(in_buffer[95]<<2)+(in_buffer[95]<<6))+(0-(in_buffer[100]<<0)-(in_buffer[100]<<2)+(in_buffer[100]<<6))+(0-(in_buffer[101]<<0)-(in_buffer[101]<<2)+(in_buffer[101]<<6))-(0-(in_buffer[107]<<0)-(in_buffer[107]<<2)+(in_buffer[107]<<6))-(0-(in_buffer[108]<<0)-(in_buffer[108]<<2)+(in_buffer[108]<<6))+(0-(in_buffer[113]<<0)-(in_buffer[113]<<2)+(in_buffer[113]<<6))-(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))+(0-(in_buffer[124]<<0)-(in_buffer[124]<<2)+(in_buffer[124]<<6))-(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6))+(0-(in_buffer[135]<<0)-(in_buffer[135]<<2)+(in_buffer[135]<<6))+(0-(in_buffer[136]<<0)-(in_buffer[136]<<2)+(in_buffer[136]<<6))+(0-(in_buffer[137]<<0)-(in_buffer[137]<<2)+(in_buffer[137]<<6))+(0-(in_buffer[140]<<0)-(in_buffer[140]<<2)+(in_buffer[140]<<6))-(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight16;
assign in_buffer_weight16=0+(0-(in_buffer[6]<<0)-(in_buffer[6]<<2)+(in_buffer[6]<<6))+(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)+(in_buffer[7]<<6))+(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)+(in_buffer[49]<<6))+(0-(in_buffer[61]<<0)-(in_buffer[61]<<2)+(in_buffer[61]<<6))+(0-(in_buffer[62]<<0)-(in_buffer[62]<<2)+(in_buffer[62]<<6))+(0-(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6))+(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)+(in_buffer[75]<<6))+(0-(in_buffer[76]<<0)-(in_buffer[76]<<2)+(in_buffer[76]<<6))+(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<2)+(in_buffer[80]<<6))+(0-(in_buffer[87]<<0)-(in_buffer[87]<<2)+(in_buffer[87]<<6))+(0-(in_buffer[88]<<0)-(in_buffer[88]<<2)+(in_buffer[88]<<6))+(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<6))+(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)+(in_buffer[90]<<6))+(0-(in_buffer[91]<<0)-(in_buffer[91]<<2)+(in_buffer[91]<<6))+(0-(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<6))-(0-(in_buffer[94]<<0)-(in_buffer[94]<<2)+(in_buffer[94]<<6))+(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6))+(0-(in_buffer[102]<<0)-(in_buffer[102]<<2)+(in_buffer[102]<<6))+(0-(in_buffer[107]<<0)-(in_buffer[107]<<2)+(in_buffer[107]<<6))+(0-(in_buffer[108]<<0)-(in_buffer[108]<<2)+(in_buffer[108]<<6))-(0-(in_buffer[113]<<0)-(in_buffer[113]<<2)+(in_buffer[113]<<6))-(0-(in_buffer[114]<<0)-(in_buffer[114]<<2)+(in_buffer[114]<<6))-(0-(in_buffer[115]<<0)-(in_buffer[115]<<2)+(in_buffer[115]<<6))-(0-(in_buffer[116]<<0)-(in_buffer[116]<<2)+(in_buffer[116]<<6))+(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))-(0-(in_buffer[124]<<0)-(in_buffer[124]<<2)+(in_buffer[124]<<6))-(0-(in_buffer[125]<<0)-(in_buffer[125]<<2)+(in_buffer[125]<<6))-(0-(in_buffer[126]<<0)-(in_buffer[126]<<2)+(in_buffer[126]<<6))-(0-(in_buffer[127]<<0)-(in_buffer[127]<<2)+(in_buffer[127]<<6))-(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))-(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight17;
assign in_buffer_weight17=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight18;
assign in_buffer_weight18=0-(0-(in_buffer[0]<<0)-(in_buffer[0]<<2)+(in_buffer[0]<<6))+(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<6))+(0-(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<6))+(0-(in_buffer[25]<<0)-(in_buffer[25]<<2)+(in_buffer[25]<<6))-(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<6))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))-(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))+(0-(in_buffer[34]<<0)-(in_buffer[34]<<2)+(in_buffer[34]<<6))+(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)+(in_buffer[36]<<6))+(0-(in_buffer[37]<<0)-(in_buffer[37]<<2)+(in_buffer[37]<<6))-(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))-(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6))+(0-(in_buffer[47]<<0)-(in_buffer[47]<<2)+(in_buffer[47]<<6))+(0-(in_buffer[48]<<0)-(in_buffer[48]<<2)+(in_buffer[48]<<6))-(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)+(in_buffer[51]<<6))+(0-(in_buffer[60]<<0)-(in_buffer[60]<<2)+(in_buffer[60]<<6))-(0-(in_buffer[62]<<0)-(in_buffer[62]<<2)+(in_buffer[62]<<6))+(0-(in_buffer[72]<<0)-(in_buffer[72]<<2)+(in_buffer[72]<<6))+(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<6))+(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight19;
assign in_buffer_weight19=0-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<6))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))-(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))+(0-(in_buffer[48]<<0)-(in_buffer[48]<<2)+(in_buffer[48]<<6))-(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))+(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight20;
assign in_buffer_weight20=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight21;
assign in_buffer_weight21=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight22;
assign in_buffer_weight22=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight23;
assign in_buffer_weight23=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight24;
assign in_buffer_weight24=0-(0-(in_buffer[26]<<0)-(in_buffer[26]<<2)+(in_buffer[26]<<6))-(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)+(in_buffer[27]<<6))-(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)+(in_buffer[38]<<6))-(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))-(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)+(in_buffer[40]<<6))-(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))-(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))-(0-(in_buffer[45]<<0)-(in_buffer[45]<<2)+(in_buffer[45]<<6))-(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))-(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)+(in_buffer[54]<<6))-(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))-(0-(in_buffer[64]<<0)-(in_buffer[64]<<2)+(in_buffer[64]<<6))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))-(0-(in_buffer[66]<<0)-(in_buffer[66]<<2)+(in_buffer[66]<<6))+(0-(in_buffer[73]<<0)-(in_buffer[73]<<2)+(in_buffer[73]<<6))+(0-(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6))+(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)+(in_buffer[75]<<6))+(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)+(in_buffer[81]<<6))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<6))-(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)+(in_buffer[84]<<6))+(0-(in_buffer[85]<<0)-(in_buffer[85]<<2)+(in_buffer[85]<<6))+(0-(in_buffer[86]<<0)-(in_buffer[86]<<2)+(in_buffer[86]<<6))+(0-(in_buffer[87]<<0)-(in_buffer[87]<<2)+(in_buffer[87]<<6))+(0-(in_buffer[88]<<0)-(in_buffer[88]<<2)+(in_buffer[88]<<6))+(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<6))+(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)+(in_buffer[90]<<6))+(0-(in_buffer[91]<<0)-(in_buffer[91]<<2)+(in_buffer[91]<<6))+(0-(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<6))+(0-(in_buffer[93]<<1)-(in_buffer[93]<<3)+(in_buffer[93]<<7))+(0-(in_buffer[94]<<0)-(in_buffer[94]<<2)+(in_buffer[94]<<6))-(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6))+(0-(in_buffer[98]<<0)-(in_buffer[98]<<2)+(in_buffer[98]<<6))+(0-(in_buffer[99]<<1)-(in_buffer[99]<<3)+(in_buffer[99]<<7))+(0-(in_buffer[100]<<1)-(in_buffer[100]<<3)+(in_buffer[100]<<7))+(0-(in_buffer[101]<<0)-(in_buffer[101]<<2)+(in_buffer[101]<<6))+(0-(in_buffer[102]<<1)-(in_buffer[102]<<3)+(in_buffer[102]<<7))+(0-(in_buffer[103]<<1)-(in_buffer[103]<<3)+(in_buffer[103]<<7))+(0-(in_buffer[104]<<0)-(in_buffer[104]<<2)+(in_buffer[104]<<6))+(0-(in_buffer[105]<<0)-(in_buffer[105]<<2)+(in_buffer[105]<<6))-(0-(in_buffer[107]<<0)-(in_buffer[107]<<2)+(in_buffer[107]<<6))+(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)+(in_buffer[112]<<6))+(0-(in_buffer[113]<<0)-(in_buffer[113]<<2)+(in_buffer[113]<<6))+(0-(in_buffer[114]<<0)-(in_buffer[114]<<2)+(in_buffer[114]<<6))+(0-(in_buffer[115]<<0)-(in_buffer[115]<<2)+(in_buffer[115]<<6))-(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<6))-(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))-(0-(in_buffer[121]<<0)-(in_buffer[121]<<2)+(in_buffer[121]<<6))-(0-(in_buffer[122]<<0)-(in_buffer[122]<<2)+(in_buffer[122]<<6))-(0-(in_buffer[123]<<0)-(in_buffer[123]<<2)+(in_buffer[123]<<6))-(0-(in_buffer[124]<<0)-(in_buffer[124]<<2)+(in_buffer[124]<<6))-(0-(in_buffer[125]<<0)-(in_buffer[125]<<2)+(in_buffer[125]<<6))-(0-(in_buffer[126]<<0)-(in_buffer[126]<<2)+(in_buffer[126]<<6))-(0-(in_buffer[127]<<0)-(in_buffer[127]<<2)+(in_buffer[127]<<6))-(0-(in_buffer[128]<<0)-(in_buffer[128]<<2)+(in_buffer[128]<<6))-(0-(in_buffer[129]<<0)-(in_buffer[129]<<2)+(in_buffer[129]<<6))-(0-(in_buffer[130]<<0)-(in_buffer[130]<<2)+(in_buffer[130]<<6))-(0-(in_buffer[136]<<0)-(in_buffer[136]<<2)+(in_buffer[136]<<6))-(0-(in_buffer[137]<<0)-(in_buffer[137]<<2)+(in_buffer[137]<<6))-(0-(in_buffer[138]<<0)-(in_buffer[138]<<2)+(in_buffer[138]<<6))-(0-(in_buffer[139]<<0)-(in_buffer[139]<<2)+(in_buffer[139]<<6))-(0-(in_buffer[140]<<0)-(in_buffer[140]<<2)+(in_buffer[140]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight25;
assign in_buffer_weight25=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight26;
assign in_buffer_weight26=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight27;
assign in_buffer_weight27=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight28;
assign in_buffer_weight28=0-(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<6))-(0-(in_buffer[16]<<0)-(in_buffer[16]<<2)+(in_buffer[16]<<6))-(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)+(in_buffer[17]<<6))-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<6))-(0-(in_buffer[21]<<0)-(in_buffer[21]<<2)+(in_buffer[21]<<6))-(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)+(in_buffer[27]<<6))-(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<6))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))-(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))-(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))-(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))-(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))-(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6))-(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))-(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))-(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))-(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)+(in_buffer[54]<<6))-(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))+(0-(in_buffer[58]<<0)-(in_buffer[58]<<2)+(in_buffer[58]<<6))+(0-(in_buffer[61]<<0)-(in_buffer[61]<<2)+(in_buffer[61]<<6))+(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)+(in_buffer[77]<<6))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6))+(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<2)+(in_buffer[80]<<6))+(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<6))-(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6))-(0-(in_buffer[107]<<0)-(in_buffer[107]<<2)+(in_buffer[107]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight29;
assign in_buffer_weight29=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight30;
assign in_buffer_weight30=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight31;
assign in_buffer_weight31=0+(0-(in_buffer[0]<<0)-(in_buffer[0]<<2)+(in_buffer[0]<<6))-(0-(in_buffer[4]<<0)-(in_buffer[4]<<2)+(in_buffer[4]<<6))-(0-(in_buffer[6]<<0)-(in_buffer[6]<<2)+(in_buffer[6]<<6))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<6))-(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<6))-(0-(in_buffer[25]<<0)-(in_buffer[25]<<2)+(in_buffer[25]<<6))+(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<6))+(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))+(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))-(0-(in_buffer[34]<<0)-(in_buffer[34]<<2)+(in_buffer[34]<<6))+(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)+(in_buffer[40]<<6))+(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))+(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))+(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6))+(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))+(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)+(in_buffer[54]<<6))+(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))+(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))-(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6))-(0-(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<6))+(0-(in_buffer[99]<<0)-(in_buffer[99]<<2)+(in_buffer[99]<<6))-(0-(in_buffer[109]<<0)-(in_buffer[109]<<2)+(in_buffer[109]<<6))+(0-(in_buffer[111]<<0)-(in_buffer[111]<<2)+(in_buffer[111]<<6))+(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)+(in_buffer[112]<<6))+(0-(in_buffer[114]<<0)-(in_buffer[114]<<2)+(in_buffer[114]<<6))+(0-(in_buffer[115]<<0)-(in_buffer[115]<<2)+(in_buffer[115]<<6))+(0-(in_buffer[116]<<0)-(in_buffer[116]<<2)+(in_buffer[116]<<6))-(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<6))-(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight32;
assign in_buffer_weight32=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight33;
assign in_buffer_weight33=0-(0-(in_buffer[0]<<0)-(in_buffer[0]<<2)+(in_buffer[0]<<6))+(0-(in_buffer[20]<<0)-(in_buffer[20]<<2)+(in_buffer[20]<<6))+(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)+(in_buffer[38]<<6))-(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))-(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))+(0-(in_buffer[61]<<0)-(in_buffer[61]<<2)+(in_buffer[61]<<6))+(0-(in_buffer[62]<<0)-(in_buffer[62]<<2)+(in_buffer[62]<<6))+(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)+(in_buffer[70]<<6))+(0-(in_buffer[71]<<0)-(in_buffer[71]<<2)+(in_buffer[71]<<6))+(0-(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight34;
assign in_buffer_weight34=0-(0-(in_buffer[8]<<0)-(in_buffer[8]<<2)+(in_buffer[8]<<6))-(0-(in_buffer[9]<<0)-(in_buffer[9]<<2)+(in_buffer[9]<<6))-(0-(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<6))-(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<6))-(0-(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<6))-(0-(in_buffer[34]<<0)-(in_buffer[34]<<2)+(in_buffer[34]<<6))-(0-(in_buffer[35]<<0)-(in_buffer[35]<<2)+(in_buffer[35]<<6))-(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)+(in_buffer[36]<<6))-(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)+(in_buffer[38]<<6))-(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)+(in_buffer[51]<<6))-(0-(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6))+(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)+(in_buffer[77]<<6))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6))+(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))+(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<6))+(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)+(in_buffer[90]<<6))+(0-(in_buffer[95]<<0)-(in_buffer[95]<<2)+(in_buffer[95]<<6))+(0-(in_buffer[107]<<0)-(in_buffer[107]<<2)+(in_buffer[107]<<6))+(0-(in_buffer[108]<<0)-(in_buffer[108]<<2)+(in_buffer[108]<<6))-(0-(in_buffer[110]<<0)-(in_buffer[110]<<2)+(in_buffer[110]<<6))-(0-(in_buffer[117]<<0)-(in_buffer[117]<<2)+(in_buffer[117]<<6))+(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))+(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<6))+(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6))+(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))+(0-(in_buffer[142]<<0)-(in_buffer[142]<<2)+(in_buffer[142]<<6))+(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight35;
assign in_buffer_weight35=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight36;
assign in_buffer_weight36=0-(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)+(in_buffer[70]<<6))-(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))-(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<6))+(0-(in_buffer[104]<<0)-(in_buffer[104]<<2)+(in_buffer[104]<<6))-(0-(in_buffer[108]<<0)-(in_buffer[108]<<2)+(in_buffer[108]<<6))-(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))-(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<6))-(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6))-(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))-(0-(in_buffer[133]<<0)-(in_buffer[133]<<2)+(in_buffer[133]<<6))-(0-(in_buffer[136]<<0)-(in_buffer[136]<<2)+(in_buffer[136]<<6))-(0-(in_buffer[137]<<0)-(in_buffer[137]<<2)+(in_buffer[137]<<6))-(0-(in_buffer[142]<<0)-(in_buffer[142]<<2)+(in_buffer[142]<<6))-(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight37;
assign in_buffer_weight37=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight38;
assign in_buffer_weight38=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight39;
assign in_buffer_weight39=0-(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))-(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))-(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)+(in_buffer[54]<<6))-(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))-(0-(in_buffer[56]<<0)-(in_buffer[56]<<2)+(in_buffer[56]<<6))-(0-(in_buffer[63]<<0)-(in_buffer[63]<<2)+(in_buffer[63]<<6))-(0-(in_buffer[64]<<0)-(in_buffer[64]<<2)+(in_buffer[64]<<6))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))-(0-(in_buffer[66]<<1)-(in_buffer[66]<<3)+(in_buffer[66]<<7))-(0-(in_buffer[67]<<0)-(in_buffer[67]<<2)+(in_buffer[67]<<6))-(0-(in_buffer[68]<<0)-(in_buffer[68]<<2)+(in_buffer[68]<<6))-(0-(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6))-(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)+(in_buffer[75]<<6))-(0-(in_buffer[76]<<0)-(in_buffer[76]<<2)+(in_buffer[76]<<6))-(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)+(in_buffer[77]<<6))-(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6))-(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))-(0-(in_buffer[80]<<0)-(in_buffer[80]<<2)+(in_buffer[80]<<6))-(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)+(in_buffer[81]<<6))+(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)+(in_buffer[84]<<6))-(0-(in_buffer[87]<<0)-(in_buffer[87]<<2)+(in_buffer[87]<<6))-(0-(in_buffer[88]<<0)-(in_buffer[88]<<2)+(in_buffer[88]<<6))-(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<6))-(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)+(in_buffer[90]<<6))-(0-(in_buffer[91]<<0)-(in_buffer[91]<<2)+(in_buffer[91]<<6))-(0-(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<6))-(0-(in_buffer[93]<<0)-(in_buffer[93]<<2)+(in_buffer[93]<<6))+(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6))-(0-(in_buffer[99]<<0)-(in_buffer[99]<<2)+(in_buffer[99]<<6))-(0-(in_buffer[101]<<0)-(in_buffer[101]<<2)+(in_buffer[101]<<6))-(0-(in_buffer[102]<<0)-(in_buffer[102]<<2)+(in_buffer[102]<<6))-(0-(in_buffer[105]<<0)-(in_buffer[105]<<2)+(in_buffer[105]<<6))+(0-(in_buffer[107]<<0)-(in_buffer[107]<<2)+(in_buffer[107]<<6))+(0-(in_buffer[108]<<0)-(in_buffer[108]<<2)+(in_buffer[108]<<6))+(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))+(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<6))+(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6))+(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))+(0-(in_buffer[133]<<0)-(in_buffer[133]<<2)+(in_buffer[133]<<6))+(0-(in_buffer[134]<<0)-(in_buffer[134]<<2)+(in_buffer[134]<<6))+(0-(in_buffer[137]<<0)-(in_buffer[137]<<2)+(in_buffer[137]<<6))+(0-(in_buffer[139]<<0)-(in_buffer[139]<<2)+(in_buffer[139]<<6))+(0-(in_buffer[140]<<0)-(in_buffer[140]<<2)+(in_buffer[140]<<6))+(0-(in_buffer[141]<<0)-(in_buffer[141]<<2)+(in_buffer[141]<<6))+(0-(in_buffer[142]<<0)-(in_buffer[142]<<2)+(in_buffer[142]<<6))+(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight40;
assign in_buffer_weight40=0+(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<6))+(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))+(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))+(0-(in_buffer[35]<<0)-(in_buffer[35]<<2)+(in_buffer[35]<<6))+(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))+(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))-(0-(in_buffer[66]<<0)-(in_buffer[66]<<2)+(in_buffer[66]<<6))+(0-(in_buffer[69]<<0)-(in_buffer[69]<<2)+(in_buffer[69]<<6))-(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6))+(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)+(in_buffer[81]<<6))+(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))+(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))+(0-(in_buffer[133]<<0)-(in_buffer[133]<<2)+(in_buffer[133]<<6))+(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight41;
assign in_buffer_weight41=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight42;
assign in_buffer_weight42=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight43;
assign in_buffer_weight43=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight44;
assign in_buffer_weight44=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight45;
assign in_buffer_weight45=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight46;
assign in_buffer_weight46=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight47;
assign in_buffer_weight47=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight48;
assign in_buffer_weight48=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight49;
assign in_buffer_weight49=0-(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<6))-(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)+(in_buffer[27]<<6))-(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<6))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))-(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))-(0-(in_buffer[31]<<0)-(in_buffer[31]<<2)+(in_buffer[31]<<6))-(0-(in_buffer[32]<<0)-(in_buffer[32]<<2)+(in_buffer[32]<<6))+(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)+(in_buffer[36]<<6))-(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))-(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)+(in_buffer[40]<<6))-(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))-(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))-(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6))-(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))-(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)+(in_buffer[51]<<6))-(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))-(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))-(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)+(in_buffer[54]<<6))-(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))-(0-(in_buffer[64]<<0)-(in_buffer[64]<<2)+(in_buffer[64]<<6))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))-(0-(in_buffer[66]<<0)-(in_buffer[66]<<2)+(in_buffer[66]<<6))-(0-(in_buffer[67]<<0)-(in_buffer[67]<<2)+(in_buffer[67]<<6))-(0-(in_buffer[68]<<0)-(in_buffer[68]<<2)+(in_buffer[68]<<6))-(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)+(in_buffer[75]<<6))-(0-(in_buffer[76]<<0)-(in_buffer[76]<<2)+(in_buffer[76]<<6))-(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)+(in_buffer[77]<<6))-(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6))-(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))-(0-(in_buffer[88]<<0)-(in_buffer[88]<<2)+(in_buffer[88]<<6))-(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<6))-(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)+(in_buffer[90]<<6))-(0-(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<6))+(0-(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<6))-(0-(in_buffer[101]<<0)-(in_buffer[101]<<2)+(in_buffer[101]<<6))-(0-(in_buffer[102]<<0)-(in_buffer[102]<<2)+(in_buffer[102]<<6))-(0-(in_buffer[115]<<0)-(in_buffer[115]<<2)+(in_buffer[115]<<6))-(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<6))-(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6))-(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))-(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight50;
assign in_buffer_weight50=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight51;
assign in_buffer_weight51=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight52;
assign in_buffer_weight52=0-(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)+(in_buffer[38]<<6))-(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<6))-(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)+(in_buffer[40]<<6))-(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))-(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)+(in_buffer[42]<<6))-(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6))-(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))-(0-(in_buffer[45]<<0)-(in_buffer[45]<<2)+(in_buffer[45]<<6))-(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)+(in_buffer[51]<<6))-(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))-(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))-(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)+(in_buffer[54]<<6))-(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))+(0-(in_buffer[58]<<0)-(in_buffer[58]<<2)+(in_buffer[58]<<6))+(0-(in_buffer[61]<<0)-(in_buffer[61]<<2)+(in_buffer[61]<<6))+(0-(in_buffer[62]<<0)-(in_buffer[62]<<2)+(in_buffer[62]<<6))+(0-(in_buffer[63]<<0)-(in_buffer[63]<<2)+(in_buffer[63]<<6))+(0-(in_buffer[64]<<0)-(in_buffer[64]<<2)+(in_buffer[64]<<6))+(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))+(0-(in_buffer[66]<<1)-(in_buffer[66]<<3)+(in_buffer[66]<<7))+(0-(in_buffer[67]<<1)-(in_buffer[67]<<3)+(in_buffer[67]<<7))+(0-(in_buffer[68]<<1)-(in_buffer[68]<<3)+(in_buffer[68]<<7))+(0-(in_buffer[69]<<0)-(in_buffer[69]<<2)+(in_buffer[69]<<6))+(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)+(in_buffer[70]<<6))+(0-(in_buffer[73]<<0)-(in_buffer[73]<<2)+(in_buffer[73]<<6))+(0-(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6))+(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)+(in_buffer[75]<<6))+(0-(in_buffer[76]<<0)-(in_buffer[76]<<2)+(in_buffer[76]<<6))+(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)+(in_buffer[77]<<6))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6))+(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<6))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<2)+(in_buffer[80]<<6))+(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)+(in_buffer[81]<<6))-(0-(in_buffer[85]<<0)-(in_buffer[85]<<2)+(in_buffer[85]<<6))-(0-(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<6))+(0-(in_buffer[128]<<0)-(in_buffer[128]<<2)+(in_buffer[128]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight53;
assign in_buffer_weight53=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight54;
assign in_buffer_weight54=0-(0-(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<6))-(0-(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<6))-(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<6))-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<6))-(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))+(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)+(in_buffer[38]<<6))+(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))+(0-(in_buffer[50]<<0)-(in_buffer[50]<<2)+(in_buffer[50]<<6))+(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)+(in_buffer[51]<<6))+(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))+(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))+(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)+(in_buffer[54]<<6))+(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<6))+(0-(in_buffer[56]<<0)-(in_buffer[56]<<2)+(in_buffer[56]<<6))+(0-(in_buffer[57]<<0)-(in_buffer[57]<<2)+(in_buffer[57]<<6))+(0-(in_buffer[64]<<0)-(in_buffer[64]<<2)+(in_buffer[64]<<6))+(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))+(0-(in_buffer[66]<<0)-(in_buffer[66]<<2)+(in_buffer[66]<<6))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<2)+(in_buffer[80]<<6))+(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)+(in_buffer[84]<<6))+(0-(in_buffer[87]<<0)-(in_buffer[87]<<2)+(in_buffer[87]<<6))+(0-(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<6))+(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6))-(0-(in_buffer[113]<<0)-(in_buffer[113]<<2)+(in_buffer[113]<<6))-(0-(in_buffer[114]<<0)-(in_buffer[114]<<2)+(in_buffer[114]<<6))-(0-(in_buffer[124]<<0)-(in_buffer[124]<<2)+(in_buffer[124]<<6))-(0-(in_buffer[125]<<0)-(in_buffer[125]<<2)+(in_buffer[125]<<6))-(0-(in_buffer[126]<<0)-(in_buffer[126]<<2)+(in_buffer[126]<<6))-(0-(in_buffer[127]<<0)-(in_buffer[127]<<2)+(in_buffer[127]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight55;
assign in_buffer_weight55=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight56;
assign in_buffer_weight56=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight57;
assign in_buffer_weight57=0+(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)+(in_buffer[27]<<6))+(0-(in_buffer[32]<<0)-(in_buffer[32]<<2)+(in_buffer[32]<<6))-(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<6))+(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<6))-(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<6))-(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<6))-(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)+(in_buffer[90]<<6))+(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)+(in_buffer[119]<<6))+(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<6))+(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6))+(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight58;
assign in_buffer_weight58=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight59;
assign in_buffer_weight59=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight60;
assign in_buffer_weight60=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight61;
assign in_buffer_weight61=0;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight62;
assign in_buffer_weight62=0+(0-(in_buffer[19]<<0)-(in_buffer[19]<<2)+(in_buffer[19]<<6))+(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<6))+(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)+(in_buffer[29]<<6))+(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<6))+(0-(in_buffer[31]<<0)-(in_buffer[31]<<2)+(in_buffer[31]<<6))+(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6))-(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<6))+(0-(in_buffer[62]<<0)-(in_buffer[62]<<2)+(in_buffer[62]<<6))-(0-(in_buffer[64]<<0)-(in_buffer[64]<<2)+(in_buffer[64]<<6))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)+(in_buffer[65]<<6))-(0-(in_buffer[66]<<0)-(in_buffer[66]<<2)+(in_buffer[66]<<6))+(0-(in_buffer[69]<<0)-(in_buffer[69]<<2)+(in_buffer[69]<<6))+(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)+(in_buffer[70]<<6))+(0-(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6))-(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)+(in_buffer[77]<<6))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<6))+(0-(in_buffer[85]<<0)-(in_buffer[85]<<2)+(in_buffer[85]<<6))+(0-(in_buffer[98]<<0)-(in_buffer[98]<<2)+(in_buffer[98]<<6))+(0-(in_buffer[105]<<0)-(in_buffer[105]<<2)+(in_buffer[105]<<6))-(0-(in_buffer[108]<<0)-(in_buffer[108]<<2)+(in_buffer[108]<<6))+(0-(in_buffer[110]<<0)-(in_buffer[110]<<2)+(in_buffer[110]<<6))+(0-(in_buffer[111]<<0)-(in_buffer[111]<<2)+(in_buffer[111]<<6))+(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)+(in_buffer[112]<<6))+(0-(in_buffer[113]<<0)-(in_buffer[113]<<2)+(in_buffer[113]<<6))+(0-(in_buffer[115]<<0)-(in_buffer[115]<<2)+(in_buffer[115]<<6))+(0-(in_buffer[116]<<0)-(in_buffer[116]<<2)+(in_buffer[116]<<6))+(0-(in_buffer[117]<<0)-(in_buffer[117]<<2)+(in_buffer[117]<<6))+(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<6))-(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<6))+(0-(in_buffer[124]<<0)-(in_buffer[124]<<2)+(in_buffer[124]<<6))+(0-(in_buffer[125]<<0)-(in_buffer[125]<<2)+(in_buffer[125]<<6))+(0-(in_buffer[127]<<0)-(in_buffer[127]<<2)+(in_buffer[127]<<6))-(0-(in_buffer[131]<<0)-(in_buffer[131]<<2)+(in_buffer[131]<<6))-(0-(in_buffer[132]<<0)-(in_buffer[132]<<2)+(in_buffer[132]<<6))-(0-(in_buffer[133]<<0)-(in_buffer[133]<<2)+(in_buffer[133]<<6))-(0-(in_buffer[134]<<0)-(in_buffer[134]<<2)+(in_buffer[134]<<6))-(0-(in_buffer[142]<<0)-(in_buffer[142]<<2)+(in_buffer[142]<<6))-(0-(in_buffer[143]<<0)-(in_buffer[143]<<2)+(in_buffer[143]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight63;
assign in_buffer_weight63=0;
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
wire signed [DATA_WIDTH-1:0]   weight_bias10;
wire signed [DATA_WIDTH-1:0]   weight_bias11;
wire signed [DATA_WIDTH-1:0]   weight_bias12;
wire signed [DATA_WIDTH-1:0]   weight_bias13;
wire signed [DATA_WIDTH-1:0]   weight_bias14;
wire signed [DATA_WIDTH-1:0]   weight_bias15;
wire signed [DATA_WIDTH-1:0]   weight_bias16;
wire signed [DATA_WIDTH-1:0]   weight_bias17;
wire signed [DATA_WIDTH-1:0]   weight_bias18;
wire signed [DATA_WIDTH-1:0]   weight_bias19;
wire signed [DATA_WIDTH-1:0]   weight_bias20;
wire signed [DATA_WIDTH-1:0]   weight_bias21;
wire signed [DATA_WIDTH-1:0]   weight_bias22;
wire signed [DATA_WIDTH-1:0]   weight_bias23;
wire signed [DATA_WIDTH-1:0]   weight_bias24;
wire signed [DATA_WIDTH-1:0]   weight_bias25;
wire signed [DATA_WIDTH-1:0]   weight_bias26;
wire signed [DATA_WIDTH-1:0]   weight_bias27;
wire signed [DATA_WIDTH-1:0]   weight_bias28;
wire signed [DATA_WIDTH-1:0]   weight_bias29;
wire signed [DATA_WIDTH-1:0]   weight_bias30;
wire signed [DATA_WIDTH-1:0]   weight_bias31;
wire signed [DATA_WIDTH-1:0]   weight_bias32;
wire signed [DATA_WIDTH-1:0]   weight_bias33;
wire signed [DATA_WIDTH-1:0]   weight_bias34;
wire signed [DATA_WIDTH-1:0]   weight_bias35;
wire signed [DATA_WIDTH-1:0]   weight_bias36;
wire signed [DATA_WIDTH-1:0]   weight_bias37;
wire signed [DATA_WIDTH-1:0]   weight_bias38;
wire signed [DATA_WIDTH-1:0]   weight_bias39;
wire signed [DATA_WIDTH-1:0]   weight_bias40;
wire signed [DATA_WIDTH-1:0]   weight_bias41;
wire signed [DATA_WIDTH-1:0]   weight_bias42;
wire signed [DATA_WIDTH-1:0]   weight_bias43;
wire signed [DATA_WIDTH-1:0]   weight_bias44;
wire signed [DATA_WIDTH-1:0]   weight_bias45;
wire signed [DATA_WIDTH-1:0]   weight_bias46;
wire signed [DATA_WIDTH-1:0]   weight_bias47;
wire signed [DATA_WIDTH-1:0]   weight_bias48;
wire signed [DATA_WIDTH-1:0]   weight_bias49;
wire signed [DATA_WIDTH-1:0]   weight_bias50;
wire signed [DATA_WIDTH-1:0]   weight_bias51;
wire signed [DATA_WIDTH-1:0]   weight_bias52;
wire signed [DATA_WIDTH-1:0]   weight_bias53;
wire signed [DATA_WIDTH-1:0]   weight_bias54;
wire signed [DATA_WIDTH-1:0]   weight_bias55;
wire signed [DATA_WIDTH-1:0]   weight_bias56;
wire signed [DATA_WIDTH-1:0]   weight_bias57;
wire signed [DATA_WIDTH-1:0]   weight_bias58;
wire signed [DATA_WIDTH-1:0]   weight_bias59;
wire signed [DATA_WIDTH-1:0]   weight_bias60;
wire signed [DATA_WIDTH-1:0]   weight_bias61;
wire signed [DATA_WIDTH-1:0]   weight_bias62;
wire signed [DATA_WIDTH-1:0]   weight_bias63;
assign weight_bias0=in_buffer_weight0+(0);
assign weight_bias1=in_buffer_weight1+(0);
assign weight_bias2=in_buffer_weight2+(0);
assign weight_bias3=in_buffer_weight3+(0);
assign weight_bias4=in_buffer_weight4+(0);
assign weight_bias5=in_buffer_weight5+(0);
assign weight_bias6=in_buffer_weight6+(-59);
assign weight_bias7=in_buffer_weight7+(0);
assign weight_bias8=in_buffer_weight8+(0);
assign weight_bias9=in_buffer_weight9+(59);
assign weight_bias10=in_buffer_weight10+(0);
assign weight_bias11=in_buffer_weight11+(0);
assign weight_bias12=in_buffer_weight12+(0);
assign weight_bias13=in_buffer_weight13+(0);
assign weight_bias14=in_buffer_weight14+(-118);
assign weight_bias15=in_buffer_weight15+(0);
assign weight_bias16=in_buffer_weight16+(59);
assign weight_bias17=in_buffer_weight17+(0);
assign weight_bias18=in_buffer_weight18+(118);
assign weight_bias19=in_buffer_weight19+(177);
assign weight_bias20=in_buffer_weight20+(0);
assign weight_bias21=in_buffer_weight21+(0);
assign weight_bias22=in_buffer_weight22+(0);
assign weight_bias23=in_buffer_weight23+(0);
assign weight_bias24=in_buffer_weight24+(0);
assign weight_bias25=in_buffer_weight25+(0);
assign weight_bias26=in_buffer_weight26+(0);
assign weight_bias27=in_buffer_weight27+(0);
assign weight_bias28=in_buffer_weight28+(118);
assign weight_bias29=in_buffer_weight29+(0);
assign weight_bias30=in_buffer_weight30+(0);
assign weight_bias31=in_buffer_weight31+(-59);
assign weight_bias32=in_buffer_weight32+(0);
assign weight_bias33=in_buffer_weight33+(-59);
assign weight_bias34=in_buffer_weight34+(118);
assign weight_bias35=in_buffer_weight35+(0);
assign weight_bias36=in_buffer_weight36+(-59);
assign weight_bias37=in_buffer_weight37+(0);
assign weight_bias38=in_buffer_weight38+(0);
assign weight_bias39=in_buffer_weight39+(-59);
assign weight_bias40=in_buffer_weight40+(59);
assign weight_bias41=in_buffer_weight41+(0);
assign weight_bias42=in_buffer_weight42+(0);
assign weight_bias43=in_buffer_weight43+(0);
assign weight_bias44=in_buffer_weight44+(0);
assign weight_bias45=in_buffer_weight45+(0);
assign weight_bias46=in_buffer_weight46+(0);
assign weight_bias47=in_buffer_weight47+(0);
assign weight_bias48=in_buffer_weight48+(0);
assign weight_bias49=in_buffer_weight49+(-59);
assign weight_bias50=in_buffer_weight50+(0);
assign weight_bias51=in_buffer_weight51+(0);
assign weight_bias52=in_buffer_weight52+(-59);
assign weight_bias53=in_buffer_weight53+(0);
assign weight_bias54=in_buffer_weight54+(-59);
assign weight_bias55=in_buffer_weight55+(0);
assign weight_bias56=in_buffer_weight56+(0);
assign weight_bias57=in_buffer_weight57+(0);
assign weight_bias58=in_buffer_weight58+(0);
assign weight_bias59=in_buffer_weight59+(0);
assign weight_bias60=in_buffer_weight60+(0);
assign weight_bias61=in_buffer_weight61+(0);
assign weight_bias62=in_buffer_weight62+(0);
assign weight_bias63=in_buffer_weight63+(0);
wire signed [DATA_WIDTH-1:0]   bias_relu0;
wire signed [DATA_WIDTH-1:0]   bias_relu1;
wire signed [DATA_WIDTH-1:0]   bias_relu2;
wire signed [DATA_WIDTH-1:0]   bias_relu3;
wire signed [DATA_WIDTH-1:0]   bias_relu4;
wire signed [DATA_WIDTH-1:0]   bias_relu5;
wire signed [DATA_WIDTH-1:0]   bias_relu6;
wire signed [DATA_WIDTH-1:0]   bias_relu7;
wire signed [DATA_WIDTH-1:0]   bias_relu8;
wire signed [DATA_WIDTH-1:0]   bias_relu9;
wire signed [DATA_WIDTH-1:0]   bias_relu10;
wire signed [DATA_WIDTH-1:0]   bias_relu11;
wire signed [DATA_WIDTH-1:0]   bias_relu12;
wire signed [DATA_WIDTH-1:0]   bias_relu13;
wire signed [DATA_WIDTH-1:0]   bias_relu14;
wire signed [DATA_WIDTH-1:0]   bias_relu15;
wire signed [DATA_WIDTH-1:0]   bias_relu16;
wire signed [DATA_WIDTH-1:0]   bias_relu17;
wire signed [DATA_WIDTH-1:0]   bias_relu18;
wire signed [DATA_WIDTH-1:0]   bias_relu19;
wire signed [DATA_WIDTH-1:0]   bias_relu20;
wire signed [DATA_WIDTH-1:0]   bias_relu21;
wire signed [DATA_WIDTH-1:0]   bias_relu22;
wire signed [DATA_WIDTH-1:0]   bias_relu23;
wire signed [DATA_WIDTH-1:0]   bias_relu24;
wire signed [DATA_WIDTH-1:0]   bias_relu25;
wire signed [DATA_WIDTH-1:0]   bias_relu26;
wire signed [DATA_WIDTH-1:0]   bias_relu27;
wire signed [DATA_WIDTH-1:0]   bias_relu28;
wire signed [DATA_WIDTH-1:0]   bias_relu29;
wire signed [DATA_WIDTH-1:0]   bias_relu30;
wire signed [DATA_WIDTH-1:0]   bias_relu31;
wire signed [DATA_WIDTH-1:0]   bias_relu32;
wire signed [DATA_WIDTH-1:0]   bias_relu33;
wire signed [DATA_WIDTH-1:0]   bias_relu34;
wire signed [DATA_WIDTH-1:0]   bias_relu35;
wire signed [DATA_WIDTH-1:0]   bias_relu36;
wire signed [DATA_WIDTH-1:0]   bias_relu37;
wire signed [DATA_WIDTH-1:0]   bias_relu38;
wire signed [DATA_WIDTH-1:0]   bias_relu39;
wire signed [DATA_WIDTH-1:0]   bias_relu40;
wire signed [DATA_WIDTH-1:0]   bias_relu41;
wire signed [DATA_WIDTH-1:0]   bias_relu42;
wire signed [DATA_WIDTH-1:0]   bias_relu43;
wire signed [DATA_WIDTH-1:0]   bias_relu44;
wire signed [DATA_WIDTH-1:0]   bias_relu45;
wire signed [DATA_WIDTH-1:0]   bias_relu46;
wire signed [DATA_WIDTH-1:0]   bias_relu47;
wire signed [DATA_WIDTH-1:0]   bias_relu48;
wire signed [DATA_WIDTH-1:0]   bias_relu49;
wire signed [DATA_WIDTH-1:0]   bias_relu50;
wire signed [DATA_WIDTH-1:0]   bias_relu51;
wire signed [DATA_WIDTH-1:0]   bias_relu52;
wire signed [DATA_WIDTH-1:0]   bias_relu53;
wire signed [DATA_WIDTH-1:0]   bias_relu54;
wire signed [DATA_WIDTH-1:0]   bias_relu55;
wire signed [DATA_WIDTH-1:0]   bias_relu56;
wire signed [DATA_WIDTH-1:0]   bias_relu57;
wire signed [DATA_WIDTH-1:0]   bias_relu58;
wire signed [DATA_WIDTH-1:0]   bias_relu59;
wire signed [DATA_WIDTH-1:0]   bias_relu60;
wire signed [DATA_WIDTH-1:0]   bias_relu61;
wire signed [DATA_WIDTH-1:0]   bias_relu62;
wire signed [DATA_WIDTH-1:0]   bias_relu63;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign bias_relu32=(weight_bias32[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias32;
assign bias_relu33=(weight_bias33[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias33;
assign bias_relu34=(weight_bias34[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias34;
assign bias_relu35=(weight_bias35[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias35;
assign bias_relu36=(weight_bias36[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias36;
assign bias_relu37=(weight_bias37[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias37;
assign bias_relu38=(weight_bias38[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias38;
assign bias_relu39=(weight_bias39[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias39;
assign bias_relu40=(weight_bias40[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias40;
assign bias_relu41=(weight_bias41[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias41;
assign bias_relu42=(weight_bias42[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias42;
assign bias_relu43=(weight_bias43[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias43;
assign bias_relu44=(weight_bias44[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias44;
assign bias_relu45=(weight_bias45[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias45;
assign bias_relu46=(weight_bias46[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias46;
assign bias_relu47=(weight_bias47[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias47;
assign bias_relu48=(weight_bias48[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias48;
assign bias_relu49=(weight_bias49[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias49;
assign bias_relu50=(weight_bias50[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias50;
assign bias_relu51=(weight_bias51[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias51;
assign bias_relu52=(weight_bias52[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias52;
assign bias_relu53=(weight_bias53[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias53;
assign bias_relu54=(weight_bias54[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias54;
assign bias_relu55=(weight_bias55[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias55;
assign bias_relu56=(weight_bias56[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias56;
assign bias_relu57=(weight_bias57[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias57;
assign bias_relu58=(weight_bias58[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias58;
assign bias_relu59=(weight_bias59[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias59;
assign bias_relu60=(weight_bias60[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias60;
assign bias_relu61=(weight_bias61[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias61;
assign bias_relu62=(weight_bias62[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias62;
assign bias_relu63=(weight_bias63[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias63;
assign layer_out={bias_relu63,bias_relu62,bias_relu61,bias_relu60,bias_relu59,bias_relu58,bias_relu57,bias_relu56,bias_relu55,bias_relu54,bias_relu53,bias_relu52,bias_relu51,bias_relu50,bias_relu49,bias_relu48,bias_relu47,bias_relu46,bias_relu45,bias_relu44,bias_relu43,bias_relu42,bias_relu41,bias_relu40,bias_relu39,bias_relu38,bias_relu37,bias_relu36,bias_relu35,bias_relu34,bias_relu33,bias_relu32,bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule