module layer2_tcb_121x32x10
(
    input clk,
    input rst,
   input valid,
   output  reg ready,
    input [25*32-1:0]  layer_in,
    output [40*10-1:0]   layer_out
);
parameter DATA_WIDTH   =   40;
reg [DATA_WIDTH-1:0]    layer_in_buffer    [0:32-1];
integer i;
always@(posedge clk )
    begin
        if(rst)
            begin
                for(i=0;i<32;i=i+1)
                    begin
                        layer_in_buffer[i]<=0;
                    end
            end
        else
        begin
       layer_in_buffer[0]<=layer_in[24:0];
       layer_in_buffer[1]<=layer_in[49:25];
       layer_in_buffer[2]<=layer_in[74:50];
       layer_in_buffer[3]<=layer_in[99:75];
       layer_in_buffer[4]<=layer_in[124:100];
       layer_in_buffer[5]<=layer_in[149:125];
       layer_in_buffer[6]<=layer_in[174:150];
       layer_in_buffer[7]<=layer_in[199:175];
       layer_in_buffer[8]<=layer_in[224:200];
       layer_in_buffer[9]<=layer_in[249:225];
       layer_in_buffer[10]<=layer_in[274:250];
       layer_in_buffer[11]<=layer_in[299:275];
       layer_in_buffer[12]<=layer_in[324:300];
       layer_in_buffer[13]<=layer_in[349:325];
       layer_in_buffer[14]<=layer_in[374:350];
       layer_in_buffer[15]<=layer_in[399:375];
       layer_in_buffer[16]<=layer_in[424:400];
       layer_in_buffer[17]<=layer_in[449:425];
       layer_in_buffer[18]<=layer_in[474:450];
       layer_in_buffer[19]<=layer_in[499:475];
       layer_in_buffer[20]<=layer_in[524:500];
       layer_in_buffer[21]<=layer_in[549:525];
       layer_in_buffer[22]<=layer_in[574:550];
       layer_in_buffer[23]<=layer_in[599:575];
       layer_in_buffer[24]<=layer_in[624:600];
       layer_in_buffer[25]<=layer_in[649:625];
       layer_in_buffer[26]<=layer_in[674:650];
       layer_in_buffer[27]<=layer_in[699:675];
       layer_in_buffer[28]<=layer_in[724:700];
       layer_in_buffer[29]<=layer_in[749:725];
       layer_in_buffer[30]<=layer_in[774:750];
       layer_in_buffer[31]<=layer_in[799:775];
        end
   end

wire [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0+(0+(layer_in_buffer[0]<<1)+(layer_in_buffer[0]<<5)-(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<11))+(0+(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<4)-(layer_in_buffer[1]<<6)-(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<12))+(0-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<6)-(layer_in_buffer[2]<<8)-(layer_in_buffer[2]<<10)+(layer_in_buffer[2]<<13))+(0+(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<7)-(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<13))+(0+(layer_in_buffer[4]<<1)+(layer_in_buffer[4]<<3)+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<10)+(layer_in_buffer[4]<<12))-(0+(layer_in_buffer[5]<<5)+(layer_in_buffer[5]<<6)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<11))-(0+(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<2)-(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<12))+(0+(layer_in_buffer[7]<<4)+(layer_in_buffer[7]<<5)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<10))-(0+(layer_in_buffer[8]<<1)+(layer_in_buffer[8]<<2)-(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<13))-(0+(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<4)-(layer_in_buffer[9]<<6)-(layer_in_buffer[9]<<9)+(layer_in_buffer[9]<<13))+(0-(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<8))-(0-(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<6)+(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<9))-(0-(layer_in_buffer[12]<<4)+(layer_in_buffer[12]<<9)+(layer_in_buffer[12]<<11)+(layer_in_buffer[12]<<12))+(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<1)-(layer_in_buffer[13]<<4)-(layer_in_buffer[13]<<6)-(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<11))-(0+(layer_in_buffer[14]<<1)+(layer_in_buffer[14]<<7)+(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<12))-(0+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<5)+(layer_in_buffer[15]<<9)+(layer_in_buffer[15]<<12))-(0+(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<3)+(layer_in_buffer[16]<<8))-(0+(layer_in_buffer[17]<<0)+(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<3)+(layer_in_buffer[17]<<9)+(layer_in_buffer[17]<<11))+(0+(layer_in_buffer[18]<<3)-(layer_in_buffer[18]<<6)+(layer_in_buffer[18]<<11))-(0+(layer_in_buffer[19]<<0)+(layer_in_buffer[19]<<1)-(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<12))-(0+(layer_in_buffer[20]<<3)+(layer_in_buffer[20]<<4)+(layer_in_buffer[20]<<7)+(layer_in_buffer[20]<<9))-(0+(layer_in_buffer[21]<<1)-(layer_in_buffer[21]<<5)-(layer_in_buffer[21]<<10)+(layer_in_buffer[21]<<13))+(0+(layer_in_buffer[22]<<1)+(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<7))-(0-(layer_in_buffer[23]<<1)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<8)+(layer_in_buffer[23]<<9))-(0+(layer_in_buffer[24]<<3)-(layer_in_buffer[24]<<6)+(layer_in_buffer[24]<<11))+(0+(layer_in_buffer[25]<<5)+(layer_in_buffer[25]<<6)+(layer_in_buffer[25]<<9)+(layer_in_buffer[25]<<11))+(0+(layer_in_buffer[26]<<1)+(layer_in_buffer[26]<<3)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<10))+(0+(layer_in_buffer[27]<<0)+(layer_in_buffer[27]<<1)-(layer_in_buffer[27]<<7)+(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<10))-(0+(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<3)-(layer_in_buffer[28]<<6)-(layer_in_buffer[28]<<8)-(layer_in_buffer[28]<<10)+(layer_in_buffer[28]<<12)+(layer_in_buffer[28]<<13))-(0+(layer_in_buffer[29]<<3)+(layer_in_buffer[29]<<4)+(layer_in_buffer[29]<<7)+(layer_in_buffer[29]<<9))-(0+(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<7)+(layer_in_buffer[30]<<14))+(0+(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<8)+(layer_in_buffer[31]<<11));
wire [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0-(0+(layer_in_buffer[0]<<1)-(layer_in_buffer[0]<<5)-(layer_in_buffer[0]<<7)+(layer_in_buffer[0]<<9)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<14))+(0-(layer_in_buffer[1]<<1)+(layer_in_buffer[1]<<6)+(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<9))+(0+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<2)-(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<10)+(layer_in_buffer[2]<<11))-(0+(layer_in_buffer[3]<<1)-(layer_in_buffer[3]<<6)+(layer_in_buffer[3]<<12)+(layer_in_buffer[3]<<14))-(0-(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<4)-(layer_in_buffer[4]<<6)-(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<11))+(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<10)+(layer_in_buffer[5]<<13))+(0-(layer_in_buffer[6]<<1)-(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<13))-(0+(layer_in_buffer[7]<<1)+(layer_in_buffer[7]<<2)-(layer_in_buffer[7]<<5)-(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<14))-(0-(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<3)+(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<10))-(0+(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<2)-(layer_in_buffer[9]<<6)+(layer_in_buffer[9]<<13))-(0-(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<3)-(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<8)+(layer_in_buffer[10]<<11))+(0+(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<10))-(0-(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<3)+(layer_in_buffer[12]<<4)-(layer_in_buffer[12]<<11)+(layer_in_buffer[12]<<14))-(0-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<9)+(layer_in_buffer[13]<<10))-(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<7)-(layer_in_buffer[14]<<9)-(layer_in_buffer[14]<<11)+(layer_in_buffer[14]<<14))+(0+(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<1)-(layer_in_buffer[15]<<4)-(layer_in_buffer[15]<<6)-(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<10)+(layer_in_buffer[15]<<11))-(0-(layer_in_buffer[16]<<1)+(layer_in_buffer[16]<<6)+(layer_in_buffer[16]<<8)+(layer_in_buffer[16]<<9))+(0-(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<10)-(layer_in_buffer[17]<<12)+(layer_in_buffer[17]<<15))-(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)-(layer_in_buffer[18]<<5)+(layer_in_buffer[18]<<8)-(layer_in_buffer[18]<<10)+(layer_in_buffer[18]<<13))-(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<7)+(layer_in_buffer[19]<<10)+(layer_in_buffer[19]<<15))+(0+(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<2)-(layer_in_buffer[20]<<4)-(layer_in_buffer[20]<<7)+(layer_in_buffer[20]<<11))-(0+(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<3)+(layer_in_buffer[21]<<6)-(layer_in_buffer[21]<<8)+(layer_in_buffer[21]<<14))-(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<4)-(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<10))+(0+(layer_in_buffer[23]<<0)+(layer_in_buffer[23]<<1)-(layer_in_buffer[23]<<7)+(layer_in_buffer[23]<<9)+(layer_in_buffer[23]<<10))+(0+(layer_in_buffer[24]<<0)+(layer_in_buffer[24]<<1)+(layer_in_buffer[24]<<4)+(layer_in_buffer[24]<<7)-(layer_in_buffer[24]<<9)+(layer_in_buffer[24]<<14))-(0-(layer_in_buffer[25]<<1)+(layer_in_buffer[25]<<5)+(layer_in_buffer[25]<<6)+(layer_in_buffer[25]<<9)+(layer_in_buffer[25]<<13))+(0+(layer_in_buffer[26]<<6)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<10)+(layer_in_buffer[26]<<12))-(0+(layer_in_buffer[27]<<0)+(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6)+(layer_in_buffer[27]<<9))-(0-(layer_in_buffer[28]<<0)-(layer_in_buffer[28]<<2)-(layer_in_buffer[28]<<4)+(layer_in_buffer[28]<<7)-(layer_in_buffer[28]<<10)+(layer_in_buffer[28]<<12)+(layer_in_buffer[28]<<13))+(0-(layer_in_buffer[29]<<0)+(layer_in_buffer[29]<<5)+(layer_in_buffer[29]<<6)-(layer_in_buffer[29]<<9)+(layer_in_buffer[29]<<11)+(layer_in_buffer[29]<<12))+(0-(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<3)+(layer_in_buffer[30]<<7)+(layer_in_buffer[30]<<11)+(layer_in_buffer[30]<<13))-(0+(layer_in_buffer[31]<<1)+(layer_in_buffer[31]<<2)-(layer_in_buffer[31]<<8)+(layer_in_buffer[31]<<10)+(layer_in_buffer[31]<<11));
wire [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0+(0+(layer_in_buffer[0]<<1)+(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<5)+(layer_in_buffer[0]<<7))-(0-(layer_in_buffer[1]<<2)-(layer_in_buffer[1]<<4)+(layer_in_buffer[1]<<9)+(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<14))-(0-(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<3)+(layer_in_buffer[2]<<5)-(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<13))-(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<7)+(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<13))+(0-(layer_in_buffer[4]<<1)+(layer_in_buffer[4]<<5)-(layer_in_buffer[4]<<7)-(layer_in_buffer[4]<<9)+(layer_in_buffer[4]<<12))-(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<3)-(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<10)+(layer_in_buffer[5]<<12)+(layer_in_buffer[5]<<13))+(0+(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<5)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<10))+(0+(layer_in_buffer[7]<<1)+(layer_in_buffer[7]<<5)-(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<11))+(0-(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<7)-(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<13))-(0+(layer_in_buffer[9]<<1)-(layer_in_buffer[9]<<4)+(layer_in_buffer[9]<<9))+(0+(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<2)-(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<8)+(layer_in_buffer[10]<<13))-(0+(layer_in_buffer[11]<<1)-(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<9))-(0+(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<4)-(layer_in_buffer[12]<<6)+(layer_in_buffer[12]<<9)+(layer_in_buffer[12]<<12))+(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<1)-(layer_in_buffer[13]<<4)-(layer_in_buffer[13]<<6)-(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<11))-(0+(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<3)-(layer_in_buffer[14]<<5)-(layer_in_buffer[14]<<8)-(layer_in_buffer[14]<<10)+(layer_in_buffer[14]<<13))+(0+(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<4)-(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<10))+(0-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<7)+(layer_in_buffer[16]<<9)+(layer_in_buffer[16]<<10))-(0-(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<3)+(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<10))+(0+(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<4)-(layer_in_buffer[18]<<7)+(layer_in_buffer[18]<<10))-(0-(layer_in_buffer[19]<<1)+(layer_in_buffer[19]<<6)+(layer_in_buffer[19]<<8)+(layer_in_buffer[19]<<9))+(0-(layer_in_buffer[20]<<1)+(layer_in_buffer[20]<<5)-(layer_in_buffer[20]<<7)-(layer_in_buffer[20]<<9)+(layer_in_buffer[20]<<12))+(0-(layer_in_buffer[21]<<0)+(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<3)+(layer_in_buffer[21]<<6)+(layer_in_buffer[21]<<8)+(layer_in_buffer[21]<<10)+(layer_in_buffer[21]<<11))-(0-(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<9)+(layer_in_buffer[22]<<10))+(0+(layer_in_buffer[23]<<2)-(layer_in_buffer[23]<<5)+(layer_in_buffer[23]<<10))+(0-(layer_in_buffer[24]<<0)-(layer_in_buffer[24]<<2)+(layer_in_buffer[24]<<5)+(layer_in_buffer[24]<<11))-(0-(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<4)+(layer_in_buffer[25]<<5)+(layer_in_buffer[25]<<8)+(layer_in_buffer[25]<<12))+(0-(layer_in_buffer[26]<<0)+(layer_in_buffer[26]<<3)-(layer_in_buffer[26]<<5)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<8)+(layer_in_buffer[26]<<11))+(0+(layer_in_buffer[27]<<0)+(layer_in_buffer[27]<<1)-(layer_in_buffer[27]<<7)+(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<10))-(0-(layer_in_buffer[28]<<1)+(layer_in_buffer[28]<<4)-(layer_in_buffer[28]<<6)+(layer_in_buffer[28]<<8)+(layer_in_buffer[28]<<9)+(layer_in_buffer[28]<<12))+(0+(layer_in_buffer[29]<<0)+(layer_in_buffer[29]<<2)-(layer_in_buffer[29]<<8)+(layer_in_buffer[29]<<11)+(layer_in_buffer[29]<<12))-(0-(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<3)+(layer_in_buffer[30]<<4)-(layer_in_buffer[30]<<11)+(layer_in_buffer[30]<<14))+(0+(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<3)+(layer_in_buffer[31]<<6)+(layer_in_buffer[31]<<8));
wire [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0-(0+(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<5)-(layer_in_buffer[0]<<7)-(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<14))-(0-(layer_in_buffer[1]<<0)+(layer_in_buffer[1]<<3)-(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<7)+(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<11))-(0-(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<3)+(layer_in_buffer[2]<<7)+(layer_in_buffer[2]<<11)+(layer_in_buffer[2]<<13))-(0+(layer_in_buffer[3]<<1)+(layer_in_buffer[3]<<2)-(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<11))-(0-(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<3)-(layer_in_buffer[4]<<5)+(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<11))+(0+(layer_in_buffer[5]<<1)-(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<7)-(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<13))+(0+(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<7)+(layer_in_buffer[6]<<9))+(0-(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<3)-(layer_in_buffer[7]<<5)+(layer_in_buffer[7]<<7)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<11))-(0+(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<3)-(layer_in_buffer[9]<<5)-(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<11))-(0+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<4)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<9)+(layer_in_buffer[10]<<11)+(layer_in_buffer[10]<<14))+(0+(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<6))+(0+(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<3)-(layer_in_buffer[12]<<9)+(layer_in_buffer[12]<<11)+(layer_in_buffer[12]<<12))+(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<4)-(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<10))-(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<3)+(layer_in_buffer[14]<<6)+(layer_in_buffer[14]<<10))+(0+(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<12))-(0+(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<3)+(layer_in_buffer[16]<<6)+(layer_in_buffer[16]<<8))-(0+(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<10)+(layer_in_buffer[17]<<13))+(0+(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<1)-(layer_in_buffer[18]<<4)-(layer_in_buffer[18]<<6)-(layer_in_buffer[18]<<8)+(layer_in_buffer[18]<<10)+(layer_in_buffer[18]<<11))-(0+(layer_in_buffer[19]<<0)+(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<4)-(layer_in_buffer[19]<<6)+(layer_in_buffer[19]<<9)+(layer_in_buffer[19]<<10)+(layer_in_buffer[19]<<14))+(0+(layer_in_buffer[20]<<3)+(layer_in_buffer[20]<<6)+(layer_in_buffer[20]<<8)+(layer_in_buffer[20]<<12)+(layer_in_buffer[20]<<13))+(0-(layer_in_buffer[21]<<0)+(layer_in_buffer[21]<<4)-(layer_in_buffer[21]<<7)-(layer_in_buffer[21]<<10)+(layer_in_buffer[21]<<13))+(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<3)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<9)+(layer_in_buffer[22]<<10))-(0+(layer_in_buffer[24]<<7)+(layer_in_buffer[24]<<8)+(layer_in_buffer[24]<<11)+(layer_in_buffer[24]<<13))-(0+(layer_in_buffer[25]<<1)+(layer_in_buffer[25]<<3)-(layer_in_buffer[25]<<9)+(layer_in_buffer[25]<<12)+(layer_in_buffer[25]<<13))+(0+(layer_in_buffer[26]<<0)+(layer_in_buffer[26]<<1)+(layer_in_buffer[26]<<4)+(layer_in_buffer[26]<<6))-(0-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<7)+(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<10))-(0+(layer_in_buffer[28]<<0)+(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<3)-(layer_in_buffer[28]<<6)-(layer_in_buffer[28]<<8)+(layer_in_buffer[28]<<13))-(0+(layer_in_buffer[29]<<1)+(layer_in_buffer[29]<<3)-(layer_in_buffer[29]<<5)-(layer_in_buffer[29]<<8)+(layer_in_buffer[29]<<12))+(0+(layer_in_buffer[30]<<1)+(layer_in_buffer[30]<<2)-(layer_in_buffer[30]<<8)+(layer_in_buffer[30]<<10)+(layer_in_buffer[30]<<11))+(0+(layer_in_buffer[31]<<2)-(layer_in_buffer[31]<<4)-(layer_in_buffer[31]<<7)+(layer_in_buffer[31]<<10)+(layer_in_buffer[31]<<12));
wire [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0+(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<8))-(0+(layer_in_buffer[1]<<1)+(layer_in_buffer[1]<<4)-(layer_in_buffer[1]<<6)-(layer_in_buffer[1]<<9)-(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<14))-(0+(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<4)-(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<11)+(layer_in_buffer[2]<<13))-(0+(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)-(layer_in_buffer[3]<<4)-(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<14))-(0+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<5)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<10))+(0-(layer_in_buffer[5]<<1)-(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<11))-(0+(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<1)-(layer_in_buffer[6]<<7)+(layer_in_buffer[6]<<9)+(layer_in_buffer[6]<<10))+(0+(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<7)+(layer_in_buffer[7]<<12))+(0-(layer_in_buffer[8]<<1)-(layer_in_buffer[8]<<3)-(layer_in_buffer[8]<<5)+(layer_in_buffer[8]<<9)+(layer_in_buffer[8]<<10))+(0-(layer_in_buffer[9]<<1)-(layer_in_buffer[9]<<3)-(layer_in_buffer[9]<<5)+(layer_in_buffer[9]<<9)+(layer_in_buffer[9]<<10))-(0-(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<3)+(layer_in_buffer[10]<<4)+(layer_in_buffer[10]<<7)-(layer_in_buffer[10]<<9)+(layer_in_buffer[10]<<12))+(0+(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<7))-(0+(layer_in_buffer[12]<<1)+(layer_in_buffer[12]<<3)+(layer_in_buffer[12]<<4)-(layer_in_buffer[12]<<7)-(layer_in_buffer[12]<<9)+(layer_in_buffer[12]<<14))-(0+(layer_in_buffer[13]<<1)-(layer_in_buffer[13]<<4)+(layer_in_buffer[13]<<9))+(0+(layer_in_buffer[14]<<1)-(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<9))+(0+(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<1)-(layer_in_buffer[15]<<5)+(layer_in_buffer[15]<<12))-(0+(layer_in_buffer[16]<<1)+(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<5)+(layer_in_buffer[16]<<7))+(0+(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<3)+(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<8))+(0+(layer_in_buffer[18]<<4)-(layer_in_buffer[18]<<7)+(layer_in_buffer[18]<<12))+(0+(layer_in_buffer[19]<<0)+(layer_in_buffer[19]<<1)+(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<7)+(layer_in_buffer[19]<<10)+(layer_in_buffer[19]<<13))-(0+(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<1)-(layer_in_buffer[20]<<4)-(layer_in_buffer[20]<<7)+(layer_in_buffer[20]<<13))+(0-(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<5)+(layer_in_buffer[21]<<11))-(0-(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<3)+(layer_in_buffer[22]<<6)+(layer_in_buffer[22]<<10))+(0+(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<3)+(layer_in_buffer[23]<<8))-(0+(layer_in_buffer[24]<<2)-(layer_in_buffer[24]<<4)-(layer_in_buffer[24]<<7)+(layer_in_buffer[24]<<10)+(layer_in_buffer[24]<<12))-(0-(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<4)+(layer_in_buffer[25]<<6)+(layer_in_buffer[25]<<12)+(layer_in_buffer[25]<<13))+(0+(layer_in_buffer[26]<<3)+(layer_in_buffer[26]<<4)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<9))+(0+(layer_in_buffer[27]<<1)-(layer_in_buffer[27]<<4)+(layer_in_buffer[27]<<9))+(0+(layer_in_buffer[28]<<1)+(layer_in_buffer[28]<<3)+(layer_in_buffer[28]<<7)+(layer_in_buffer[28]<<10))+(0-(layer_in_buffer[29]<<1)-(layer_in_buffer[29]<<3)-(layer_in_buffer[29]<<5)+(layer_in_buffer[29]<<9)+(layer_in_buffer[29]<<10))+(0-(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<3)+(layer_in_buffer[30]<<4)+(layer_in_buffer[30]<<7)-(layer_in_buffer[30]<<9)+(layer_in_buffer[30]<<12))+(0+(layer_in_buffer[31]<<0)+(layer_in_buffer[31]<<1)+(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0+(0+(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<5)+(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<9)+(layer_in_buffer[0]<<12))-(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<5)-(layer_in_buffer[1]<<8)-(layer_in_buffer[1]<<10)+(layer_in_buffer[1]<<13)+(layer_in_buffer[1]<<14))+(0+(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<11))+(0-(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)-(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<9))-(0+(layer_in_buffer[4]<<1)+(layer_in_buffer[4]<<3)+(layer_in_buffer[4]<<4)-(layer_in_buffer[4]<<7)-(layer_in_buffer[4]<<9)+(layer_in_buffer[4]<<14))+(0+(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<5)+(layer_in_buffer[5]<<8)+(layer_in_buffer[5]<<10))+(0-(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<11))+(0+(layer_in_buffer[7]<<1)-(layer_in_buffer[7]<<4)-(layer_in_buffer[7]<<7)-(layer_in_buffer[7]<<10)+(layer_in_buffer[7]<<12)+(layer_in_buffer[7]<<13))+(0-(layer_in_buffer[8]<<1)+(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<9))-(0+(layer_in_buffer[9]<<0)+(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<5)+(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<11))+(0+(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<2)-(layer_in_buffer[10]<<4)-(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<11))-(0+(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<4)-(layer_in_buffer[11]<<7)+(layer_in_buffer[11]<<10))+(0+(layer_in_buffer[12]<<1)+(layer_in_buffer[12]<<3)-(layer_in_buffer[12]<<5)-(layer_in_buffer[12]<<8)+(layer_in_buffer[12]<<12))-(0+(layer_in_buffer[13]<<3)+(layer_in_buffer[13]<<5)-(layer_in_buffer[13]<<7)-(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<14))+(0+(layer_in_buffer[14]<<2)-(layer_in_buffer[14]<<5)+(layer_in_buffer[14]<<10))-(0-(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<13))-(0+(layer_in_buffer[16]<<0)+(layer_in_buffer[16]<<1)-(layer_in_buffer[16]<<7)+(layer_in_buffer[16]<<9)+(layer_in_buffer[16]<<10))+(0+(layer_in_buffer[17]<<0)+(layer_in_buffer[17]<<3)+(layer_in_buffer[17]<<4)+(layer_in_buffer[17]<<7)+(layer_in_buffer[17]<<8)+(layer_in_buffer[17]<<11)+(layer_in_buffer[17]<<14))-(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<5)+(layer_in_buffer[18]<<14))+(0+(layer_in_buffer[19]<<0)+(layer_in_buffer[19]<<1)+(layer_in_buffer[19]<<4)+(layer_in_buffer[19]<<6))+(0+(layer_in_buffer[20]<<0)-(layer_in_buffer[20]<<3)+(layer_in_buffer[20]<<5)+(layer_in_buffer[20]<<6)-(layer_in_buffer[20]<<9)+(layer_in_buffer[20]<<13)+(layer_in_buffer[20]<<14))-(0+(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<3)+(layer_in_buffer[21]<<6)+(layer_in_buffer[21]<<8))-(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<4)-(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<10))-(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<3)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<10))+(0-(layer_in_buffer[24]<<1)-(layer_in_buffer[24]<<4)+(layer_in_buffer[24]<<9)+(layer_in_buffer[24]<<12)+(layer_in_buffer[24]<<13))+(0-(layer_in_buffer[25]<<2)-(layer_in_buffer[25]<<4)+(layer_in_buffer[25]<<7)+(layer_in_buffer[25]<<13))-(0-(layer_in_buffer[26]<<2)+(layer_in_buffer[26]<<6)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<10)+(layer_in_buffer[26]<<14))-(0-(layer_in_buffer[27]<<0)+(layer_in_buffer[27]<<5)+(layer_in_buffer[27]<<7)+(layer_in_buffer[27]<<8))+(0-(layer_in_buffer[28]<<0)+(layer_in_buffer[28]<<4)-(layer_in_buffer[28]<<7)-(layer_in_buffer[28]<<10)+(layer_in_buffer[28]<<13))-(0-(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<5)-(layer_in_buffer[29]<<8)+(layer_in_buffer[29]<<12)+(layer_in_buffer[29]<<14))-(0-(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<3)-(layer_in_buffer[30]<<6)+(layer_in_buffer[30]<<10)+(layer_in_buffer[30]<<12))+(0-(layer_in_buffer[31]<<0)+(layer_in_buffer[31]<<3)+(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<7)+(layer_in_buffer[31]<<8)+(layer_in_buffer[31]<<13)+(layer_in_buffer[31]<<14));
wire [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0+(0-(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<6)+(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<11))+(0+(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<4)-(layer_in_buffer[1]<<6)-(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<12))-(0-(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<3)+(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<10)+(layer_in_buffer[2]<<11))+(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<3)+(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<13))+(0+(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<5)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<10))-(0-(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<13))-(0+(layer_in_buffer[6]<<1)+(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<12))+(0+(layer_in_buffer[7]<<1)+(layer_in_buffer[7]<<2)-(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<10)+(layer_in_buffer[7]<<11))-(0+(layer_in_buffer[8]<<3)+(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<7)-(layer_in_buffer[8]<<9)-(layer_in_buffer[8]<<11)+(layer_in_buffer[8]<<13)+(layer_in_buffer[8]<<14))+(0-(layer_in_buffer[9]<<1)-(layer_in_buffer[9]<<3)-(layer_in_buffer[9]<<5)+(layer_in_buffer[9]<<9)+(layer_in_buffer[9]<<10))-(0+(layer_in_buffer[10]<<2)-(layer_in_buffer[10]<<4)-(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<12))-(0+(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<4)-(layer_in_buffer[11]<<7)+(layer_in_buffer[11]<<10))+(0-(layer_in_buffer[12]<<2)-(layer_in_buffer[12]<<4)-(layer_in_buffer[12]<<6)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<11))+(0+(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<4)+(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<11))+(0+(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<1)-(layer_in_buffer[14]<<7)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<10))+(0-(layer_in_buffer[15]<<1)-(layer_in_buffer[15]<<4)+(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<11))-(0+(layer_in_buffer[16]<<0)+(layer_in_buffer[16]<<1)+(layer_in_buffer[16]<<4)+(layer_in_buffer[16]<<6))-(0+(layer_in_buffer[17]<<1)+(layer_in_buffer[17]<<4)+(layer_in_buffer[17]<<8)+(layer_in_buffer[17]<<13))+(0+(layer_in_buffer[18]<<5)+(layer_in_buffer[18]<<6)+(layer_in_buffer[18]<<9)+(layer_in_buffer[18]<<11))-(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<4)+(layer_in_buffer[19]<<7)-(layer_in_buffer[19]<<10)+(layer_in_buffer[19]<<12)+(layer_in_buffer[19]<<13))-(0+(layer_in_buffer[20]<<1)+(layer_in_buffer[20]<<4)-(layer_in_buffer[20]<<6)-(layer_in_buffer[20]<<9)-(layer_in_buffer[20]<<11)+(layer_in_buffer[20]<<14))-(0+(layer_in_buffer[21]<<5)-(layer_in_buffer[21]<<8)+(layer_in_buffer[21]<<13))+(0+(layer_in_buffer[22]<<1)+(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<7))+(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<3)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<10))+(0+(layer_in_buffer[24]<<1)+(layer_in_buffer[24]<<2)-(layer_in_buffer[24]<<8)+(layer_in_buffer[24]<<10)+(layer_in_buffer[24]<<11))-(0+(layer_in_buffer[25]<<0)-(layer_in_buffer[25]<<4)-(layer_in_buffer[25]<<6)+(layer_in_buffer[25]<<8)+(layer_in_buffer[25]<<9)+(layer_in_buffer[25]<<13))-(0+(layer_in_buffer[26]<<1)+(layer_in_buffer[26]<<3)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<10))+(0+(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<2)-(layer_in_buffer[27]<<5)+(layer_in_buffer[27]<<8)+(layer_in_buffer[27]<<10))+(0-(layer_in_buffer[28]<<1)-(layer_in_buffer[28]<<3)-(layer_in_buffer[28]<<5)-(layer_in_buffer[28]<<7)+(layer_in_buffer[28]<<12)+(layer_in_buffer[28]<<13))+(0-(layer_in_buffer[29]<<1)-(layer_in_buffer[29]<<3)-(layer_in_buffer[29]<<5)+(layer_in_buffer[29]<<9)+(layer_in_buffer[29]<<10))-(0+(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<2)-(layer_in_buffer[30]<<4)-(layer_in_buffer[30]<<6)+(layer_in_buffer[30]<<9)+(layer_in_buffer[30]<<10)+(layer_in_buffer[30]<<14))-(0-(layer_in_buffer[31]<<0)+(layer_in_buffer[31]<<4)-(layer_in_buffer[31]<<6)-(layer_in_buffer[31]<<8)+(layer_in_buffer[31]<<11));
wire [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0-(0-(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<6)+(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<11))-(0-(layer_in_buffer[1]<<0)+(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<6)+(layer_in_buffer[1]<<12)+(layer_in_buffer[1]<<15))+(0+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<2)-(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<10)+(layer_in_buffer[2]<<11))+(0+(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6)-(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<12))-(0+(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<6)+(layer_in_buffer[4]<<11)+(layer_in_buffer[4]<<12))+(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<5)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<10))-(0+(layer_in_buffer[6]<<0)-(layer_in_buffer[6]<<4)-(layer_in_buffer[6]<<9)+(layer_in_buffer[6]<<12))-(0-(layer_in_buffer[7]<<1)-(layer_in_buffer[7]<<5)-(layer_in_buffer[7]<<7)-(layer_in_buffer[7]<<9)-(layer_in_buffer[7]<<11)+(layer_in_buffer[7]<<15))+(0+(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<1)-(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<6)-(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<11))+(0+(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<12))+(0+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<3)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<10))-(0-(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<6)+(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<9))+(0+(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<3)+(layer_in_buffer[12]<<9)+(layer_in_buffer[12]<<11))+(0-(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<4)+(layer_in_buffer[13]<<5)+(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<12))+(0+(layer_in_buffer[14]<<1)+(layer_in_buffer[14]<<5)-(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<11))-(0+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<12)+(layer_in_buffer[15]<<13))-(0+(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<3)+(layer_in_buffer[16]<<8))-(0+(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<7)+(layer_in_buffer[17]<<10)+(layer_in_buffer[17]<<12))-(0+(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<3)-(layer_in_buffer[18]<<6)-(layer_in_buffer[18]<<9)+(layer_in_buffer[18]<<11)+(layer_in_buffer[18]<<12))+(0-(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<8)+(layer_in_buffer[19]<<12))-(0-(layer_in_buffer[20]<<1)+(layer_in_buffer[20]<<4)+(layer_in_buffer[20]<<6)-(layer_in_buffer[20]<<10)+(layer_in_buffer[20]<<14))+(0-(layer_in_buffer[21]<<0)+(layer_in_buffer[21]<<3)+(layer_in_buffer[21]<<4)+(layer_in_buffer[21]<<7)-(layer_in_buffer[21]<<9)+(layer_in_buffer[21]<<12))+(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<3)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<9)+(layer_in_buffer[22]<<10))+(0+(layer_in_buffer[23]<<0)+(layer_in_buffer[23]<<3)+(layer_in_buffer[23]<<5)+(layer_in_buffer[23]<<9)+(layer_in_buffer[23]<<10))-(0-(layer_in_buffer[24]<<3)-(layer_in_buffer[24]<<5)+(layer_in_buffer[24]<<8)+(layer_in_buffer[24]<<14))+(0-(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<3)+(layer_in_buffer[25]<<5)-(layer_in_buffer[25]<<9)+(layer_in_buffer[25]<<13))-(0+(layer_in_buffer[26]<<0)+(layer_in_buffer[26]<<3)+(layer_in_buffer[26]<<4)+(layer_in_buffer[26]<<13))-(0+(layer_in_buffer[27]<<3)+(layer_in_buffer[27]<<4)+(layer_in_buffer[27]<<7)+(layer_in_buffer[27]<<9))-(0+(layer_in_buffer[28]<<2)+(layer_in_buffer[28]<<8)+(layer_in_buffer[28]<<9)+(layer_in_buffer[28]<<13))+(0+(layer_in_buffer[29]<<0)+(layer_in_buffer[29]<<2)-(layer_in_buffer[29]<<4)-(layer_in_buffer[29]<<6)+(layer_in_buffer[29]<<9)+(layer_in_buffer[29]<<10)+(layer_in_buffer[29]<<14))+(0+(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<5)+(layer_in_buffer[30]<<7)+(layer_in_buffer[30]<<11)+(layer_in_buffer[30]<<12))-(0+(layer_in_buffer[31]<<1)-(layer_in_buffer[31]<<3)+(layer_in_buffer[31]<<7)+(layer_in_buffer[31]<<8)-(layer_in_buffer[31]<<12)+(layer_in_buffer[31]<<15));
wire [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0+(0+(layer_in_buffer[0]<<1)+(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<6)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<11))-(0+(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<7)+(layer_in_buffer[1]<<9)+(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<13))+(0+(layer_in_buffer[2]<<3)-(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<11))+(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<1)-(layer_in_buffer[3]<<4)-(layer_in_buffer[3]<<6)-(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<11))+(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<5)+(layer_in_buffer[4]<<8)-(layer_in_buffer[4]<<10)+(layer_in_buffer[4]<<13))-(0+(layer_in_buffer[5]<<1)+(layer_in_buffer[5]<<2)-(layer_in_buffer[5]<<5)-(layer_in_buffer[5]<<7)-(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<11)+(layer_in_buffer[5]<<12))-(0+(layer_in_buffer[6]<<1)+(layer_in_buffer[6]<<2)-(layer_in_buffer[6]<<9)+(layer_in_buffer[6]<<13)+(layer_in_buffer[6]<<14))-(0+(layer_in_buffer[7]<<2)-(layer_in_buffer[7]<<5)+(layer_in_buffer[7]<<10))+(0+(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<5)+(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<10)-(layer_in_buffer[8]<<12)+(layer_in_buffer[8]<<15))+(0-(layer_in_buffer[9]<<2)-(layer_in_buffer[9]<<4)-(layer_in_buffer[9]<<6)+(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<11))-(0-(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<4)-(layer_in_buffer[10]<<7)-(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<13))-(0+(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<6))+(0+(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<3)+(layer_in_buffer[12]<<8))-(0-(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<5)-(layer_in_buffer[13]<<8)-(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<12)+(layer_in_buffer[13]<<13))+(0+(layer_in_buffer[14]<<1)+(layer_in_buffer[14]<<2)-(layer_in_buffer[14]<<5)-(layer_in_buffer[14]<<7)-(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<11)+(layer_in_buffer[14]<<12))+(0+(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<11))-(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)-(layer_in_buffer[16]<<4)+(layer_in_buffer[16]<<8)+(layer_in_buffer[16]<<9))+(0-(layer_in_buffer[17]<<3)-(layer_in_buffer[17]<<5)-(layer_in_buffer[17]<<7)+(layer_in_buffer[17]<<11)+(layer_in_buffer[17]<<12))-(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)-(layer_in_buffer[18]<<4)+(layer_in_buffer[18]<<8)+(layer_in_buffer[18]<<9))+(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<3)+(layer_in_buffer[19]<<8)+(layer_in_buffer[19]<<11)+(layer_in_buffer[19]<<12))+(0+(layer_in_buffer[20]<<1)+(layer_in_buffer[20]<<3)+(layer_in_buffer[20]<<6)+(layer_in_buffer[20]<<8)+(layer_in_buffer[20]<<11)+(layer_in_buffer[20]<<12))+(0+(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<6)-(layer_in_buffer[21]<<9)+(layer_in_buffer[21]<<12))+(0-(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<8))-(0+(layer_in_buffer[23]<<1)+(layer_in_buffer[23]<<3)+(layer_in_buffer[23]<<7)+(layer_in_buffer[23]<<10))-(0+(layer_in_buffer[24]<<0)+(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<5)+(layer_in_buffer[24]<<9)+(layer_in_buffer[24]<<10))-(0+(layer_in_buffer[25]<<1)+(layer_in_buffer[25]<<7)+(layer_in_buffer[25]<<8)+(layer_in_buffer[25]<<12))+(0-(layer_in_buffer[26]<<0)+(layer_in_buffer[26]<<4)+(layer_in_buffer[26]<<5)+(layer_in_buffer[26]<<8)+(layer_in_buffer[26]<<12))+(0+(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<3)+(layer_in_buffer[27]<<8))-(0+(layer_in_buffer[28]<<0)+(layer_in_buffer[28]<<3)+(layer_in_buffer[28]<<6)-(layer_in_buffer[28]<<11)+(layer_in_buffer[28]<<15))-(0+(layer_in_buffer[29]<<0)+(layer_in_buffer[29]<<2)-(layer_in_buffer[29]<<4)+(layer_in_buffer[29]<<8)+(layer_in_buffer[29]<<12)+(layer_in_buffer[29]<<13))-(0+(layer_in_buffer[30]<<5)+(layer_in_buffer[30]<<6)+(layer_in_buffer[30]<<9)+(layer_in_buffer[30]<<11))-(0-(layer_in_buffer[31]<<3)+(layer_in_buffer[31]<<7)-(layer_in_buffer[31]<<9)-(layer_in_buffer[31]<<11)+(layer_in_buffer[31]<<14));
wire [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0+(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<8))-(0-(layer_in_buffer[1]<<1)+(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<6)+(layer_in_buffer[1]<<9)+(layer_in_buffer[1]<<13))+(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<7)+(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<12))-(0-(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)-(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<7)-(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<12)+(layer_in_buffer[3]<<13))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<5)+(layer_in_buffer[4]<<11))+(0-(layer_in_buffer[5]<<3)-(layer_in_buffer[5]<<5)-(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<11)+(layer_in_buffer[5]<<12))-(0+(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<5)+(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<12)+(layer_in_buffer[6]<<14))-(0+(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<5)+(layer_in_buffer[7]<<7)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<15))-(0-(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<3)-(layer_in_buffer[8]<<7)+(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<11)+(layer_in_buffer[8]<<14))-(0+(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<3)+(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<10))+(0+(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<4)+(layer_in_buffer[10]<<5)-(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<13))-(0+(layer_in_buffer[11]<<3)+(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<7)+(layer_in_buffer[11]<<9))+(0-(layer_in_buffer[12]<<1)-(layer_in_buffer[12]<<4)+(layer_in_buffer[12]<<7)+(layer_in_buffer[12]<<11))+(0-(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<3)+(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<11))+(0-(layer_in_buffer[14]<<3)+(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<10)+(layer_in_buffer[14]<<11))-(0-(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<3)-(layer_in_buffer[15]<<5)+(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<11))+(0+(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<3)+(layer_in_buffer[16]<<8))-(0+(layer_in_buffer[17]<<1)+(layer_in_buffer[17]<<4)+(layer_in_buffer[17]<<10)-(layer_in_buffer[17]<<12)+(layer_in_buffer[17]<<15))-(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<6)+(layer_in_buffer[18]<<7)+(layer_in_buffer[18]<<12)+(layer_in_buffer[18]<<14))+(0+(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<3)-(layer_in_buffer[19]<<9)+(layer_in_buffer[19]<<11)+(layer_in_buffer[19]<<12))-(0+(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<3)+(layer_in_buffer[20]<<6)+(layer_in_buffer[20]<<8)+(layer_in_buffer[20]<<10)+(layer_in_buffer[20]<<13))+(0+(layer_in_buffer[21]<<1)+(layer_in_buffer[21]<<3)-(layer_in_buffer[21]<<5)-(layer_in_buffer[21]<<8)+(layer_in_buffer[21]<<12))-(0+(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<3)+(layer_in_buffer[22]<<6)+(layer_in_buffer[22]<<8))-(0+(layer_in_buffer[23]<<0)+(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<9))-(0+(layer_in_buffer[24]<<0)-(layer_in_buffer[24]<<2)-(layer_in_buffer[24]<<5)+(layer_in_buffer[24]<<8)+(layer_in_buffer[24]<<10))-(0-(layer_in_buffer[25]<<0)-(layer_in_buffer[25]<<3)+(layer_in_buffer[25]<<8)+(layer_in_buffer[25]<<11)+(layer_in_buffer[25]<<12))-(0+(layer_in_buffer[26]<<4)+(layer_in_buffer[26]<<5)+(layer_in_buffer[26]<<8)+(layer_in_buffer[26]<<10))+(0-(layer_in_buffer[27]<<0)-(layer_in_buffer[27]<<3)+(layer_in_buffer[27]<<6)+(layer_in_buffer[27]<<10))+(0-(layer_in_buffer[28]<<3)-(layer_in_buffer[28]<<5)-(layer_in_buffer[28]<<7)+(layer_in_buffer[28]<<11)+(layer_in_buffer[28]<<12))-(0-(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<5)-(layer_in_buffer[29]<<8)+(layer_in_buffer[29]<<12)+(layer_in_buffer[29]<<14))+(0+(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<2)-(layer_in_buffer[30]<<5)+(layer_in_buffer[30]<<7)+(layer_in_buffer[30]<<8)+(layer_in_buffer[30]<<13))-(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<2)-(layer_in_buffer[31]<<4)-(layer_in_buffer[31]<<6)+(layer_in_buffer[31]<<11)+(layer_in_buffer[31]<<12));
wire [DATA_WIDTH-1:0]   weight_bias0;
assign weight_bias0=in_buffer_weight0+(4731);
wire [DATA_WIDTH-1:0]   weight_bias1;
assign weight_bias1=in_buffer_weight1+(747);
wire [DATA_WIDTH-1:0]   weight_bias2;
assign weight_bias2=in_buffer_weight2+(-830);
wire [DATA_WIDTH-1:0]   weight_bias3;
assign weight_bias3=in_buffer_weight3+(3901);
wire [DATA_WIDTH-1:0]   weight_bias4;
assign weight_bias4=in_buffer_weight4+(-6142);
wire [DATA_WIDTH-1:0]   weight_bias5;
assign weight_bias5=in_buffer_weight5+(1826);
wire [DATA_WIDTH-1:0]   weight_bias6;
assign weight_bias6=in_buffer_weight6+(-498);
wire [DATA_WIDTH-1:0]   weight_bias7;
assign weight_bias7=in_buffer_weight7+(4316);
wire [DATA_WIDTH-1:0]   weight_bias8;
assign weight_bias8=in_buffer_weight8+(2573);
wire [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias9=in_buffer_weight9+(-4316);
assign layer_out={
            weight_bias9,
            weight_bias8,
            weight_bias7,
            weight_bias6,
            weight_bias5,
            weight_bias4,
            weight_bias3,
            weight_bias2,
            weight_bias1,
            weight_bias0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule
