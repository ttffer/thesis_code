`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/22/2022 03:54:19 PM
// Design Name: 
// Module Name: n37sys4x4_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module n37sys4x4_testbench(

    );
    reg [17:0] word0,word1,word2,word3,word4,word5,word6,word7,word8,word9,word10,word11,word12,word13,word14,word15;
    wire [12:0]d_word0,d_word1,d_word2,d_word3,d_word4,d_word5,d_word6,d_word7,d_word8,d_word9,d_word10,d_word11,d_word12,d_word13,d_word14,d_word15;
    
    n37sys_4x4 DUT_n37(.IN0(word0),.IN1(word1),.IN2(word2),.IN3(word3),.IN4(word4),.IN5(word5),.IN6(word6),.IN7(word7),.IN8(word8),.IN9(word9),.IN10(word10),.IN11(word11),.IN12(word12),.IN13(word13),.IN14(word14),.IN15(word15),.OUT0(d_word0),.OUT1(d_word1),.OUT2(d_word2),.OUT3(d_word3),.OUT4(d_word4),.OUT5(d_word5),.OUT6(d_word6),.OUT7(d_word7),.OUT8(d_word8),.OUT9(d_word9),.OUT10(d_word10),.OUT11(d_word11),.OUT12(d_word12),.OUT13(d_word13),.OUT14(d_word14),.OUT15(d_word15));
    
    
    initial begin 
    //possible codeword
    word0='d37;word1='d37;word2='d37;word3='d37;word4='d37;word5='d37;word6='d37;word7='d37;word8='d37;word9='d37;word10='d37;word11='d37;word12='d37;word13='d37;word14='d37;word15='d37;
    #10 word0='d37;
#10 word0='d74;
#10 word0='d111;
#10 word0='d148;
#10 word0='d185;
#10 word0='d222;
#10 word0='d259;
#10 word0='d296;
#10 word0='d333;
#10 word0='d370;
#10 word0='d407;
#10 word0='d444;
#10 word0='d481;
#10 word0='d518;
#10 word0='d555;
#10 word0='d592;
#10 word0='d629;
#10 word0='d666;
#10 word0='d703;
#10 word0='d740;
#10 word0='d777;
#10 word0='d814;
#10 word0='d851;
#10 word0='d888;
#10 word0='d925;
#10 word0='d962;
#10 word0='d999;
#10 word0='d1036;
#10 word0='d1073;
#10 word0='d1110;
#10 word0='d1147;
#10 word0='d1184;
#10 word0='d1221;
#10 word0='d1258;
#10 word0='d1295;
#10 word0='d1332;
#10 word0='d1369;
#10 word0='d1406;
#10 word0='d1443;
#10 word0='d1480;
#10 word0='d1517;
#10 word0='d1554;
#10 word0='d1591;
#10 word0='d1628;
#10 word0='d1665;
#10 word0='d1702;
#10 word0='d1739;
#10 word0='d1776;
#10 word0='d1813;
#10 word0='d1850;
#10 word0='d1887;
#10 word0='d1924;
#10 word0='d1961;
#10 word0='d1998;
#10 word0='d2035;
#10 word0='d2072;
#10 word0='d2109;
#10 word0='d2146;
#10 word0='d2183;
#10 word0='d2220;
#10 word0='d2257;
#10 word0='d2294;
#10 word0='d2331;
#10 word0='d2368;
#10 word0='d2405;
#10 word0='d2442;
#10 word0='d2479;
#10 word0='d2516;
#10 word0='d2553;
#10 word0='d2590;
#10 word0='d2627;
#10 word0='d2664;
#10 word0='d2701;
#10 word0='d2738;
#10 word0='d2775;
#10 word0='d2812;
#10 word0='d2849;
#10 word0='d2886;
#10 word0='d2923;
#10 word0='d2960;
#10 word0='d2997;
#10 word0='d3034;
#10 word0='d3071;
#10 word0='d3108;
#10 word0='d3145;
#10 word0='d3182;
#10 word0='d3219;
#10 word0='d3256;
#10 word0='d3293;
#10 word0='d3330;
#10 word0='d3367;
#10 word0='d3404;
#10 word0='d3441;
#10 word0='d3478;
#10 word0='d3515;
#10 word0='d3552;
#10 word0='d3589;
#10 word0='d3626;
#10 word0='d3663;
#10 word0='d3700;
#10 word0='d3737;
#10 word0='d3774;
#10 word0='d3811;
#10 word0='d3848;
#10 word0='d3885;
#10 word0='d3922;
#10 word0='d3959;
#10 word0='d3996;
#10 word0='d4033;
#10 word0='d4070;
#10 word0='d4107;
#10 word0='d4144;
#10 word0='d4181;
#10 word0='d4218;
#10 word0='d4255;
#10 word0='d4292;
#10 word0='d4329;
#10 word0='d4366;
#10 word0='d4403;
#10 word0='d4440;
#10 word0='d4477;
#10 word0='d4514;
#10 word0='d4551;
#10 word0='d4588;
#10 word0='d4625;
#10 word0='d4662;
#10 word0='d4699;
#10 word0='d4736;
#10 word0='d4773;
#10 word0='d4810;
#10 word0='d4847;
#10 word0='d4884;
#10 word0='d4921;
#10 word0='d4958;
#10 word0='d4995;
#10 word0='d5032;
#10 word0='d5069;
#10 word0='d5106;
#10 word0='d5143;
#10 word0='d5180;
#10 word0='d5217;
#10 word0='d5254;
#10 word0='d5291;
#10 word0='d5328;
#10 word0='d5365;
#10 word0='d5402;
#10 word0='d5439;
#10 word0='d5476;
#10 word0='d5513;
#10 word0='d5550;
#10 word0='d5587;
#10 word0='d5624;
#10 word0='d5661;
#10 word0='d5698;
#10 word0='d5735;
#10 word0='d5772;
#10 word0='d5809;
#10 word0='d5846;
#10 word0='d5883;
#10 word0='d5920;
#10 word0='d5957;
#10 word0='d5994;
#10 word0='d6031;
#10 word0='d6068;
#10 word0='d6105;
#10 word0='d6142;
#10 word0='d6179;
#10 word0='d6216;
#10 word0='d6253;
#10 word0='d6290;
#10 word0='d6327;
#10 word0='d6364;
#10 word0='d6401;
#10 word0='d6438;
#10 word0='d6475;
#10 word0='d6512;
#10 word0='d6549;
#10 word0='d6586;
#10 word0='d6623;
#10 word0='d6660;
#10 word0='d6697;
#10 word0='d6734;
#10 word0='d6771;
#10 word0='d6808;
#10 word0='d6845;
#10 word0='d6882;
#10 word0='d6919;
#10 word0='d6956;
#10 word0='d6993;
#10 word0='d7030;
#10 word0='d7067;
#10 word0='d7104;
#10 word0='d7141;
#10 word0='d7178;
#10 word0='d7215;
#10 word0='d7252;
#10 word0='d7289;
#10 word0='d7326;
#10 word0='d7363;
#10 word0='d7400;
#10 word0='d7437;
#10 word0='d7474;
#10 word0='d7511;
#10 word0='d7548;
#10 word0='d7585;
#10 word0='d7622;
#10 word0='d7659;
#10 word0='d7696;
#10 word0='d7733;
#10 word0='d7770;
#10 word0='d7807;
#10 word0='d7844;
#10 word0='d7881;
#10 word0='d7918;
#10 word0='d7955;
#10 word0='d7992;
#10 word0='d8029;
#10 word0='d8066;
#10 word0='d8103;
#10 word0='d8140;
#10 word0='d8177;
#10 word0='d8214;
#10 word0='d8251;
#10 word0='d8288;
#10 word0='d8325;
#10 word0='d8362;
#10 word0='d8399;
#10 word0='d8436;
#10 word0='d8473;
#10 word0='d8510;
#10 word0='d8547;
#10 word0='d8584;
#10 word0='d8621;
#10 word0='d8658;
#10 word0='d8695;
#10 word0='d8732;
#10 word0='d8769;
#10 word0='d8806;
#10 word0='d8843;
#10 word0='d8880;
#10 word0='d8917;
#10 word0='d8954;
#10 word0='d8991;
#10 word0='d9028;
#10 word0='d9065;
#10 word0='d9102;
#10 word0='d9139;
#10 word0='d9176;
#10 word0='d9213;
#10 word0='d9250;
#10 word0='d9287;
#10 word0='d9324;
#10 word0='d9361;
#10 word0='d9398;
#10 word0='d9435;
#10 word0='d9472;
#10 word0='d9509;
#10 word0='d9546;
#10 word0='d9583;
#10 word0='d9620;
#10 word0='d9657;
#10 word0='d9694;
#10 word0='d9731;
#10 word0='d9768;
#10 word0='d9805;
#10 word0='d9842;
#10 word0='d9879;
#10 word0='d9916;
#10 word0='d9953;
#10 word0='d9990;
#10 word0='d10027;
#10 word0='d10064;
#10 word0='d10101;
#10 word0='d10138;
#10 word0='d10175;
#10 word0='d10212;
#10 word0='d10249;
#10 word0='d10286;
#10 word0='d10323;
#10 word0='d10360;
#10 word0='d10397;
#10 word0='d10434;
#10 word0='d10471;
#10 word0='d10508;
#10 word0='d10545;
#10 word0='d10582;
#10 word0='d10619;
#10 word0='d10656;
#10 word0='d10693;
#10 word0='d10730;
#10 word0='d10767;
#10 word0='d10804;
#10 word0='d10841;
#10 word0='d10878;
#10 word0='d10915;
#10 word0='d10952;
#10 word0='d10989;
#10 word0='d11026;
#10 word0='d11063;
#10 word0='d11100;
#10 word0='d11137;
#10 word0='d11174;
#10 word0='d11211;
#10 word0='d11248;
#10 word0='d11285;
#10 word0='d11322;
#10 word0='d11359;
#10 word0='d11396;
#10 word0='d11433;
#10 word0='d11470;
#10 word0='d11507;
#10 word0='d11544;
#10 word0='d11581;
#10 word0='d11618;
#10 word0='d11655;
#10 word0='d11692;
#10 word0='d11729;
#10 word0='d11766;
#10 word0='d11803;
#10 word0='d11840;
#10 word0='d11877;
#10 word0='d11914;
#10 word0='d11951;
#10 word0='d11988;
#10 word0='d12025;
#10 word0='d12062;
#10 word0='d12099;
#10 word0='d12136;
#10 word0='d12173;
#10 word0='d12210;
#10 word0='d12247;
#10 word0='d12284;
#10 word0='d12321;
#10 word0='d12358;
#10 word0='d12395;
#10 word0='d12432;
#10 word0='d12469;
#10 word0='d12506;
#10 word0='d12543;
#10 word0='d12580;
#10 word0='d12617;
#10 word0='d12654;
#10 word0='d12691;
#10 word0='d12728;
#10 word0='d12765;
#10 word0='d12802;
#10 word0='d12839;
#10 word0='d12876;
#10 word0='d12913;
#10 word0='d12950;
#10 word0='d12987;
#10 word0='d13024;
#10 word0='d13061;
#10 word0='d13098;
#10 word0='d13135;
#10 word0='d13172;
#10 word0='d13209;
#10 word0='d13246;
#10 word0='d13283;
#10 word0='d13320;
#10 word0='d13357;
#10 word0='d13394;
#10 word0='d13431;
#10 word0='d13468;
#10 word0='d13505;
#10 word0='d13542;
#10 word0='d13579;
#10 word0='d13616;
#10 word0='d13653;
#10 word0='d13690;
#10 word0='d13727;
#10 word0='d13764;
#10 word0='d13801;
#10 word0='d13838;
#10 word0='d13875;
#10 word0='d13912;
#10 word0='d13949;
#10 word0='d13986;
#10 word0='d14023;
#10 word0='d14060;
#10 word0='d14097;
#10 word0='d14134;
#10 word0='d14171;
#10 word0='d14208;
#10 word0='d14245;
#10 word0='d14282;
#10 word0='d14319;
#10 word0='d14356;
#10 word0='d14393;
#10 word0='d14430;
#10 word0='d14467;
#10 word0='d14504;
#10 word0='d14541;
#10 word0='d14578;
#10 word0='d14615;
#10 word0='d14652;
#10 word0='d14689;
#10 word0='d14726;
#10 word0='d14763;
#10 word0='d14800;
#10 word0='d14837;
#10 word0='d14874;
#10 word0='d14911;
#10 word0='d14948;
#10 word0='d14985;
#10 word0='d15022;
#10 word0='d15059;
#10 word0='d15096;
#10 word0='d15133;
#10 word0='d15170;
#10 word0='d15207;
#10 word0='d15244;
#10 word0='d15281;
#10 word0='d15318;
#10 word0='d15355;
#10 word0='d15392;
#10 word0='d15429;
#10 word0='d15466;
#10 word0='d15503;
#10 word0='d15540;
#10 word0='d15577;
#10 word0='d15614;
#10 word0='d15651;
#10 word0='d15688;
#10 word0='d15725;
#10 word0='d15762;
#10 word0='d15799;
#10 word0='d15836;
#10 word0='d15873;
#10 word0='d15910;
#10 word0='d15947;
#10 word0='d15984;
#10 word0='d16021;
#10 word0='d16058;
#10 word0='d16095;
#10 word0='d16132;
#10 word0='d16169;
#10 word0='d16206;
#10 word0='d16243;
#10 word0='d16280;
#10 word0='d16317;
#10 word0='d16354;
#10 word0='d16391;
#10 word0='d16428;
#10 word0='d16465;
#10 word0='d16502;
#10 word0='d16539;
#10 word0='d16576;
#10 word0='d16613;
#10 word0='d16650;
#10 word0='d16687;
#10 word0='d16724;
#10 word0='d16761;
#10 word0='d16798;
#10 word0='d16835;
#10 word0='d16872;
#10 word0='d16909;
#10 word0='d16946;
#10 word0='d16983;
#10 word0='d17020;
#10 word0='d17057;
#10 word0='d17094;
#10 word0='d17131;
#10 word0='d17168;
#10 word0='d17205;
#10 word0='d17242;
#10 word0='d17279;
#10 word0='d17316;
#10 word0='d17353;
#10 word0='d17390;
#10 word0='d17427;
#10 word0='d17464;
#10 word0='d17501;
#10 word0='d17538;
#10 word0='d17575;
#10 word0='d17612;
#10 word0='d17649;
#10 word0='d17686;
#10 word0='d17723;
#10 word0='d17760;
#10 word0='d17797;
#10 word0='d17834;
#10 word0='d17871;
#10 word0='d17908;
#10 word0='d17945;
#10 word0='d17982;
#10 word0='d18019;
#10 word0='d18056;
#10 word0='d18093;
#10 word0='d18130;
#10 word0='d18167;
#10 word0='d18204;
#10 word0='d18241;
#10 word0='d18278;
#10 word0='d18315;
#10 word0='d18352;
#10 word0='d18389;
#10 word0='d18426;
#10 word0='d18463;
#10 word0='d18500;
#10 word0='d18537;
#10 word0='d18574;
#10 word0='d18611;
#10 word0='d18648;
#10 word0='d18685;
#10 word0='d18722;
#10 word0='d18759;
#10 word0='d18796;
#10 word0='d18833;
#10 word0='d18870;
#10 word0='d18907;
#10 word0='d18944;
#10 word0='d18981;
#10 word0='d19018;
#10 word0='d19055;
#10 word0='d19092;
#10 word0='d19129;
#10 word0='d19166;
#10 word0='d19203;
#10 word0='d19240;
#10 word0='d19277;
#10 word0='d19314;
#10 word0='d19351;
#10 word0='d19388;
#10 word0='d19425;
#10 word0='d19462;
#10 word0='d19499;
#10 word0='d19536;
#10 word0='d19573;
#10 word0='d19610;
#10 word0='d19647;
#10 word0='d19684;
#10 word0='d19721;
#10 word0='d19758;
#10 word0='d19795;
#10 word0='d19832;
#10 word0='d19869;
#10 word0='d19906;
#10 word0='d19943;
#10 word0='d19980;
#10 word0='d20017;
#10 word0='d20054;
#10 word0='d20091;
#10 word0='d20128;
#10 word0='d20165;
#10 word0='d20202;
#10 word0='d20239;
#10 word0='d20276;
#10 word0='d20313;
#10 word0='d20350;
#10 word0='d20387;
#10 word0='d20424;
#10 word0='d20461;
#10 word0='d20498;
#10 word0='d20535;
#10 word0='d20572;
#10 word0='d20609;
#10 word0='d20646;
#10 word0='d20683;
#10 word0='d20720;
#10 word0='d20757;
#10 word0='d20794;
#10 word0='d20831;
#10 word0='d20868;
#10 word0='d20905;
#10 word0='d20942;
#10 word0='d20979;
#10 word0='d21016;
#10 word0='d21053;
#10 word0='d21090;
#10 word0='d21127;
#10 word0='d21164;
#10 word0='d21201;
#10 word0='d21238;
#10 word0='d21275;
#10 word0='d21312;
#10 word0='d21349;
#10 word0='d21386;
#10 word0='d21423;
#10 word0='d21460;
#10 word0='d21497;
#10 word0='d21534;
#10 word0='d21571;
#10 word0='d21608;
#10 word0='d21645;
#10 word0='d21682;
#10 word0='d21719;
#10 word0='d21756;
#10 word0='d21793;
#10 word0='d21830;
#10 word0='d21867;
#10 word0='d21904;
#10 word0='d21941;
#10 word0='d21978;
#10 word0='d22015;
#10 word0='d22052;
#10 word0='d22089;
#10 word0='d22126;
#10 word0='d22163;
#10 word0='d22200;
#10 word0='d22237;
#10 word0='d22274;
#10 word0='d22311;
#10 word0='d22348;
#10 word0='d22385;
#10 word0='d22422;
#10 word0='d22459;
#10 word0='d22496;
#10 word0='d22533;
#10 word0='d22570;
#10 word0='d22607;
#10 word0='d22644;
#10 word0='d22681;
#10 word0='d22718;
#10 word0='d22755;
#10 word0='d22792;
#10 word0='d22829;
#10 word0='d22866;
#10 word0='d22903;
#10 word0='d22940;
#10 word0='d22977;
#10 word0='d23014;
#10 word0='d23051;
#10 word0='d23088;
#10 word0='d23125;
#10 word0='d23162;
#10 word0='d23199;
#10 word0='d23236;
#10 word0='d23273;
#10 word0='d23310;
#10 word0='d23347;
#10 word0='d23384;
#10 word0='d23421;
#10 word0='d23458;
#10 word0='d23495;
#10 word0='d23532;
#10 word0='d23569;
#10 word0='d23606;
#10 word0='d23643;
#10 word0='d23680;
#10 word0='d23717;
#10 word0='d23754;
#10 word0='d23791;
#10 word0='d23828;
#10 word0='d23865;
#10 word0='d23902;
#10 word0='d23939;
#10 word0='d23976;
#10 word0='d24013;
#10 word0='d24050;
#10 word0='d24087;
#10 word0='d24124;
#10 word0='d24161;
#10 word0='d24198;
#10 word0='d24235;
#10 word0='d24272;
#10 word0='d24309;
#10 word0='d24346;
#10 word0='d24383;
#10 word0='d24420;
#10 word0='d24457;
#10 word0='d24494;
#10 word0='d24531;
#10 word0='d24568;
#10 word0='d24605;
#10 word0='d24642;
#10 word0='d24679;
#10 word0='d24716;
#10 word0='d24753;
#10 word0='d24790;
#10 word0='d24827;
#10 word0='d24864;
#10 word0='d24901;
#10 word0='d24938;
#10 word0='d24975;
#10 word0='d25012;
#10 word0='d25049;
#10 word0='d25086;
#10 word0='d25123;
#10 word0='d25160;
#10 word0='d25197;
#10 word0='d25234;
#10 word0='d25271;
#10 word0='d25308;
#10 word0='d25345;
#10 word0='d25382;
#10 word0='d25419;
#10 word0='d25456;
#10 word0='d25493;
#10 word0='d25530;
#10 word0='d25567;
#10 word0='d25604;
#10 word0='d25641;
#10 word0='d25678;
#10 word0='d25715;
#10 word0='d25752;
#10 word0='d25789;
#10 word0='d25826;
#10 word0='d25863;
#10 word0='d25900;
#10 word0='d25937;
#10 word0='d25974;
#10 word0='d26011;
#10 word0='d26048;
#10 word0='d26085;
#10 word0='d26122;
#10 word0='d26159;
#10 word0='d26196;
#10 word0='d26233;
#10 word0='d26270;
#10 word0='d26307;
#10 word0='d26344;
#10 word0='d26381;
#10 word0='d26418;
#10 word0='d26455;
#10 word0='d26492;
#10 word0='d26529;
#10 word0='d26566;
#10 word0='d26603;
#10 word0='d26640;
#10 word0='d26677;
#10 word0='d26714;
#10 word0='d26751;
#10 word0='d26788;
#10 word0='d26825;
#10 word0='d26862;
#10 word0='d26899;
#10 word0='d26936;
#10 word0='d26973;
#10 word0='d27010;
#10 word0='d27047;
#10 word0='d27084;
#10 word0='d27121;
#10 word0='d27158;
#10 word0='d27195;
#10 word0='d27232;
#10 word0='d27269;
#10 word0='d27306;
#10 word0='d27343;
#10 word0='d27380;
#10 word0='d27417;
#10 word0='d27454;
#10 word0='d27491;
#10 word0='d27528;
#10 word0='d27565;
#10 word0='d27602;
#10 word0='d27639;
#10 word0='d27676;
#10 word0='d27713;
#10 word0='d27750;
#10 word0='d27787;
#10 word0='d27824;
#10 word0='d27861;
#10 word0='d27898;
#10 word0='d27935;
#10 word0='d27972;
#10 word0='d28009;
#10 word0='d28046;
#10 word0='d28083;
#10 word0='d28120;
#10 word0='d28157;
#10 word0='d28194;
#10 word0='d28231;
#10 word0='d28268;
#10 word0='d28305;
#10 word0='d28342;
#10 word0='d28379;
#10 word0='d28416;
#10 word0='d28453;
#10 word0='d28490;
#10 word0='d28527;
#10 word0='d28564;
#10 word0='d28601;
#10 word0='d28638;
#10 word0='d28675;
#10 word0='d28712;
#10 word0='d28749;
#10 word0='d28786;
#10 word0='d28823;
#10 word0='d28860;
#10 word0='d28897;
#10 word0='d28934;
#10 word0='d28971;
#10 word0='d29008;
#10 word0='d29045;
#10 word0='d29082;
#10 word0='d29119;
#10 word0='d29156;
#10 word0='d29193;
#10 word0='d29230;
#10 word0='d29267;
#10 word0='d29304;
#10 word0='d29341;
#10 word0='d29378;
#10 word0='d29415;
#10 word0='d29452;
#10 word0='d29489;
#10 word0='d29526;
#10 word0='d29563;
#10 word0='d29600;
#10 word0='d29637;
#10 word0='d29674;
#10 word0='d29711;
#10 word0='d29748;
#10 word0='d29785;
#10 word0='d29822;
#10 word0='d29859;
#10 word0='d29896;
#10 word0='d29933;
#10 word0='d29970;
#10 word0='d30007;
#10 word0='d30044;
#10 word0='d30081;
#10 word0='d30118;
#10 word0='d30155;
#10 word0='d30192;
#10 word0='d30229;
#10 word0='d30266;
#10 word0='d30303;
#10 word0='d30340;
#10 word0='d30377;
#10 word0='d30414;
#10 word0='d30451;
#10 word0='d30488;
#10 word0='d30525;
#10 word0='d30562;
#10 word0='d30599;
#10 word0='d30636;
#10 word0='d30673;
#10 word0='d30710;
#10 word0='d30747;
#10 word0='d30784;
#10 word0='d30821;
#10 word0='d30858;
#10 word0='d30895;
#10 word0='d30932;
#10 word0='d30969;
#10 word0='d31006;
#10 word0='d31043;
#10 word0='d31080;
#10 word0='d31117;
#10 word0='d31154;
#10 word0='d31191;
#10 word0='d31228;
#10 word0='d31265;
#10 word0='d31302;
#10 word0='d31339;
#10 word0='d31376;
#10 word0='d31413;
#10 word0='d31450;
#10 word0='d31487;
#10 word0='d31524;
#10 word0='d31561;
#10 word0='d31598;
#10 word0='d31635;
#10 word0='d31672;
#10 word0='d31709;
#10 word0='d31746;
#10 word0='d31783;
#10 word0='d31820;
#10 word0='d31857;
#10 word0='d31894;
#10 word0='d31931;
#10 word0='d31968;
#10 word0='d32005;
#10 word0='d32042;
#10 word0='d32079;
#10 word0='d32116;
#10 word0='d32153;
#10 word0='d32190;
#10 word0='d32227;
#10 word0='d32264;
#10 word0='d32301;
#10 word0='d32338;
#10 word0='d32375;
#10 word0='d32412;
#10 word0='d32449;
#10 word0='d32486;
#10 word0='d32523;
#10 word0='d32560;
#10 word0='d32597;
#10 word0='d32634;
#10 word0='d32671;
#10 word0='d32708;
#10 word0='d32745;
#10 word0='d32782;
#10 word0='d32819;
#10 word0='d32856;
#10 word0='d32893;
#10 word0='d32930;
#10 word0='d32967;
#10 word0='d33004;
#10 word0='d33041;
#10 word0='d33078;
#10 word0='d33115;
#10 word0='d33152;
#10 word0='d33189;
#10 word0='d33226;
#10 word0='d33263;
#10 word0='d33300;
#10 word0='d33337;
#10 word0='d33374;
#10 word0='d33411;
#10 word0='d33448;
#10 word0='d33485;
#10 word0='d33522;
#10 word0='d33559;
#10 word0='d33596;
#10 word0='d33633;
#10 word0='d33670;
#10 word0='d33707;
#10 word0='d33744;
#10 word0='d33781;
#10 word0='d33818;
#10 word0='d33855;
#10 word0='d33892;
#10 word0='d33929;
#10 word0='d33966;
#10 word0='d34003;
#10 word0='d34040;
#10 word0='d34077;
#10 word0='d34114;
#10 word0='d34151;
#10 word0='d34188;
#10 word0='d34225;
#10 word0='d34262;
#10 word0='d34299;
#10 word0='d34336;
#10 word0='d34373;
#10 word0='d34410;
#10 word0='d34447;
#10 word0='d34484;
#10 word0='d34521;
#10 word0='d34558;
#10 word0='d34595;
#10 word0='d34632;
#10 word0='d34669;
#10 word0='d34706;
#10 word0='d34743;
#10 word0='d34780;
#10 word0='d34817;
#10 word0='d34854;
#10 word0='d34891;
#10 word0='d34928;
#10 word0='d34965;
#10 word0='d35002;
#10 word0='d35039;
#10 word0='d35076;
#10 word0='d35113;
#10 word0='d35150;
#10 word0='d35187;
#10 word0='d35224;
#10 word0='d35261;
#10 word0='d35298;
#10 word0='d35335;
#10 word0='d35372;
#10 word0='d35409;
#10 word0='d35446;
#10 word0='d35483;
#10 word0='d35520;
#10 word0='d35557;
#10 word0='d35594;
#10 word0='d35631;
#10 word0='d35668;
#10 word0='d35705;
#10 word0='d35742;
#10 word0='d35779;
#10 word0='d35816;
#10 word0='d35853;
#10 word0='d35890;
#10 word0='d35927;
#10 word0='d35964;
#10 word0='d36001;
#10 word0='d36038;
#10 word0='d36075;
#10 word0='d36112;
#10 word0='d36149;
#10 word0='d36186;
#10 word0='d36223;
#10 word0='d36260;
#10 word0='d36297;
#10 word0='d36334;
#10 word0='d36371;
#10 word0='d36408;
#10 word0='d36445;
#10 word0='d36482;
#10 word0='d36519;
#10 word0='d36556;
#10 word0='d36593;
#10 word0='d36630;
#10 word0='d36667;
#10 word0='d36704;
#10 word0='d36741;
#10 word0='d36778;
#10 word0='d36815;
#10 word0='d36852;
#10 word0='d36889;
#10 word0='d36926;
#10 word0='d36963;
#10 word0='d37000;
#10 word0='d37037;
#10 word0='d37074;
#10 word0='d37111;
#10 word0='d37148;
#10 word0='d37185;
#10 word0='d37222;
#10 word0='d37259;
#10 word0='d37296;
#10 word0='d37333;
#10 word0='d37370;
#10 word0='d37407;
#10 word0='d37444;
#10 word0='d37481;
#10 word0='d37518;
#10 word0='d37555;
#10 word0='d37592;
#10 word0='d37629;
#10 word0='d37666;
#10 word0='d37703;
#10 word0='d37740;
#10 word0='d37777;
#10 word0='d37814;
#10 word0='d37851;
#10 word0='d37888;
#10 word0='d37925;
#10 word0='d37962;
#10 word0='d37999;
#10 word0='d38036;
#10 word0='d38073;
#10 word0='d38110;
#10 word0='d38147;
#10 word0='d38184;
#10 word0='d38221;
#10 word0='d38258;
#10 word0='d38295;
#10 word0='d38332;
#10 word0='d38369;
#10 word0='d38406;
#10 word0='d38443;
#10 word0='d38480;
#10 word0='d38517;
#10 word0='d38554;
#10 word0='d38591;
#10 word0='d38628;
#10 word0='d38665;
#10 word0='d38702;
#10 word0='d38739;
#10 word0='d38776;
#10 word0='d38813;
#10 word0='d38850;
#10 word0='d38887;
#10 word0='d38924;
#10 word0='d38961;
#10 word0='d38998;
#10 word0='d39035;
#10 word0='d39072;
#10 word0='d39109;
#10 word0='d39146;
#10 word0='d39183;
#10 word0='d39220;
#10 word0='d39257;
#10 word0='d39294;
#10 word0='d39331;
#10 word0='d39368;
#10 word0='d39405;
#10 word0='d39442;
#10 word0='d39479;
#10 word0='d39516;
#10 word0='d39553;
#10 word0='d39590;
#10 word0='d39627;
#10 word0='d39664;
#10 word0='d39701;
#10 word0='d39738;
#10 word0='d39775;
#10 word0='d39812;
#10 word0='d39849;
#10 word0='d39886;
#10 word0='d39923;
#10 word0='d39960;
#10 word0='d39997;
#10 word0='d40034;
#10 word0='d40071;
#10 word0='d40108;
#10 word0='d40145;
#10 word0='d40182;
#10 word0='d40219;
#10 word0='d40256;
#10 word0='d40293;
#10 word0='d40330;
#10 word0='d40367;
#10 word0='d40404;
#10 word0='d40441;
#10 word0='d40478;
#10 word0='d40515;
#10 word0='d40552;
#10 word0='d40589;
#10 word0='d40626;
#10 word0='d40663;
#10 word0='d40700;
#10 word0='d40737;
#10 word0='d40774;
#10 word0='d40811;
#10 word0='d40848;
#10 word0='d40885;
#10 word0='d40922;
#10 word0='d40959;
#10 word0='d40996;
#10 word0='d41033;
#10 word0='d41070;
#10 word0='d41107;
#10 word0='d41144;
#10 word0='d41181;
#10 word0='d41218;
#10 word0='d41255;
#10 word0='d41292;
#10 word0='d41329;
#10 word0='d41366;
#10 word0='d41403;
#10 word0='d41440;
#10 word0='d41477;
#10 word0='d41514;
#10 word0='d41551;
#10 word0='d41588;
#10 word0='d41625;
#10 word0='d41662;
#10 word0='d41699;
#10 word0='d41736;
#10 word0='d41773;
#10 word0='d41810;
#10 word0='d41847;
#10 word0='d41884;
#10 word0='d41921;
#10 word0='d41958;
#10 word0='d41995;
#10 word0='d42032;
#10 word0='d42069;
#10 word0='d42106;
#10 word0='d42143;
#10 word0='d42180;
#10 word0='d42217;
#10 word0='d42254;
#10 word0='d42291;
#10 word0='d42328;
#10 word0='d42365;
#10 word0='d42402;
#10 word0='d42439;
#10 word0='d42476;
#10 word0='d42513;
#10 word0='d42550;
#10 word0='d42587;
#10 word0='d42624;
#10 word0='d42661;
#10 word0='d42698;
#10 word0='d42735;
#10 word0='d42772;
#10 word0='d42809;
#10 word0='d42846;
#10 word0='d42883;
#10 word0='d42920;
#10 word0='d42957;
#10 word0='d42994;
#10 word0='d43031;
#10 word0='d43068;
#10 word0='d43105;
#10 word0='d43142;
#10 word0='d43179;
#10 word0='d43216;
#10 word0='d43253;
#10 word0='d43290;
#10 word0='d43327;
#10 word0='d43364;
#10 word0='d43401;
#10 word0='d43438;
#10 word0='d43475;
#10 word0='d43512;
#10 word0='d43549;
#10 word0='d43586;
#10 word0='d43623;
#10 word0='d43660;
#10 word0='d43697;
#10 word0='d43734;
#10 word0='d43771;
#10 word0='d43808;
#10 word0='d43845;
#10 word0='d43882;
#10 word0='d43919;
#10 word0='d43956;
#10 word0='d43993;
#10 word0='d44030;
#10 word0='d44067;
#10 word0='d44104;
#10 word0='d44141;
#10 word0='d44178;
#10 word0='d44215;
#10 word0='d44252;
#10 word0='d44289;
#10 word0='d44326;
#10 word0='d44363;
#10 word0='d44400;
#10 word0='d44437;
#10 word0='d44474;
#10 word0='d44511;
#10 word0='d44548;
#10 word0='d44585;
#10 word0='d44622;
#10 word0='d44659;
#10 word0='d44696;
#10 word0='d44733;
#10 word0='d44770;
#10 word0='d44807;
#10 word0='d44844;
#10 word0='d44881;
#10 word0='d44918;
#10 word0='d44955;
#10 word0='d44992;
#10 word0='d45029;
#10 word0='d45066;
#10 word0='d45103;
#10 word0='d45140;
#10 word0='d45177;
#10 word0='d45214;
#10 word0='d45251;
#10 word0='d45288;
#10 word0='d45325;
#10 word0='d45362;
#10 word0='d45399;
#10 word0='d45436;
#10 word0='d45473;
#10 word0='d45510;
#10 word0='d45547;
#10 word0='d45584;
#10 word0='d45621;
#10 word0='d45658;
#10 word0='d45695;
#10 word0='d45732;
#10 word0='d45769;
#10 word0='d45806;
#10 word0='d45843;
#10 word0='d45880;
#10 word0='d45917;
#10 word0='d45954;
#10 word0='d45991;
#10 word0='d46028;
#10 word0='d46065;
#10 word0='d46102;
#10 word0='d46139;
#10 word0='d46176;
#10 word0='d46213;
#10 word0='d46250;
#10 word0='d46287;
#10 word0='d46324;
#10 word0='d46361;
#10 word0='d46398;
#10 word0='d46435;
#10 word0='d46472;
#10 word0='d46509;
#10 word0='d46546;
#10 word0='d46583;
#10 word0='d46620;
#10 word0='d46657;
#10 word0='d46694;
#10 word0='d46731;
#10 word0='d46768;
#10 word0='d46805;
#10 word0='d46842;
#10 word0='d46879;
#10 word0='d46916;
#10 word0='d46953;
#10 word0='d46990;
#10 word0='d47027;
#10 word0='d47064;
#10 word0='d47101;
#10 word0='d47138;
#10 word0='d47175;
#10 word0='d47212;
#10 word0='d47249;
#10 word0='d47286;
#10 word0='d47323;
#10 word0='d47360;
#10 word0='d47397;
#10 word0='d47434;
#10 word0='d47471;
#10 word0='d47508;
#10 word0='d47545;
#10 word0='d47582;
#10 word0='d47619;
#10 word0='d47656;
#10 word0='d47693;
#10 word0='d47730;
#10 word0='d47767;
#10 word0='d47804;
#10 word0='d47841;
#10 word0='d47878;
#10 word0='d47915;
#10 word0='d47952;
#10 word0='d47989;
#10 word0='d48026;
#10 word0='d48063;
#10 word0='d48100;
#10 word0='d48137;
#10 word0='d48174;
#10 word0='d48211;
#10 word0='d48248;
#10 word0='d48285;
#10 word0='d48322;
#10 word0='d48359;
#10 word0='d48396;
#10 word0='d48433;
#10 word0='d48470;
#10 word0='d48507;
#10 word0='d48544;
#10 word0='d48581;
#10 word0='d48618;
#10 word0='d48655;
#10 word0='d48692;
#10 word0='d48729;
#10 word0='d48766;
#10 word0='d48803;
#10 word0='d48840;
#10 word0='d48877;
#10 word0='d48914;
#10 word0='d48951;
#10 word0='d48988;
#10 word0='d49025;
#10 word0='d49062;
#10 word0='d49099;
#10 word0='d49136;
#10 word0='d49173;
#10 word0='d49210;
#10 word0='d49247;
#10 word0='d49284;
#10 word0='d49321;
#10 word0='d49358;
#10 word0='d49395;
#10 word0='d49432;
#10 word0='d49469;
#10 word0='d49506;
#10 word0='d49543;
#10 word0='d49580;
#10 word0='d49617;
#10 word0='d49654;
#10 word0='d49691;
#10 word0='d49728;
#10 word0='d49765;
#10 word0='d49802;
#10 word0='d49839;
#10 word0='d49876;
#10 word0='d49913;
#10 word0='d49950;
#10 word0='d49987;
#10 word0='d50024;
#10 word0='d50061;
#10 word0='d50098;
#10 word0='d50135;
#10 word0='d50172;
#10 word0='d50209;
#10 word0='d50246;
#10 word0='d50283;
#10 word0='d50320;
#10 word0='d50357;
#10 word0='d50394;
#10 word0='d50431;
#10 word0='d50468;
#10 word0='d50505;
#10 word0='d50542;
#10 word0='d50579;
#10 word0='d50616;
#10 word0='d50653;
#10 word0='d50690;
#10 word0='d50727;
#10 word0='d50764;
#10 word0='d50801;
#10 word0='d50838;
#10 word0='d50875;
#10 word0='d50912;
#10 word0='d50949;
#10 word0='d50986;
#10 word0='d51023;
#10 word0='d51060;
#10 word0='d51097;
#10 word0='d51134;
#10 word0='d51171;
#10 word0='d51208;
#10 word0='d51245;
#10 word0='d51282;
#10 word0='d51319;
#10 word0='d51356;
#10 word0='d51393;
#10 word0='d51430;
#10 word0='d51467;
#10 word0='d51504;
#10 word0='d51541;
#10 word0='d51578;
#10 word0='d51615;
#10 word0='d51652;
#10 word0='d51689;
#10 word0='d51726;
#10 word0='d51763;
#10 word0='d51800;
#10 word0='d51837;
#10 word0='d51874;
#10 word0='d51911;
#10 word0='d51948;
#10 word0='d51985;
#10 word0='d52022;
#10 word0='d52059;
#10 word0='d52096;
#10 word0='d52133;
#10 word0='d52170;
#10 word0='d52207;
#10 word0='d52244;
#10 word0='d52281;
#10 word0='d52318;
#10 word0='d52355;
#10 word0='d52392;
#10 word0='d52429;
#10 word0='d52466;
#10 word0='d52503;
#10 word0='d52540;
#10 word0='d52577;
#10 word0='d52614;
#10 word0='d52651;
#10 word0='d52688;
#10 word0='d52725;
#10 word0='d52762;
#10 word0='d52799;
#10 word0='d52836;
#10 word0='d52873;
#10 word0='d52910;
#10 word0='d52947;
#10 word0='d52984;
#10 word0='d53021;
#10 word0='d53058;
#10 word0='d53095;
#10 word0='d53132;
#10 word0='d53169;
#10 word0='d53206;
#10 word0='d53243;
#10 word0='d53280;
#10 word0='d53317;
#10 word0='d53354;
#10 word0='d53391;
#10 word0='d53428;
#10 word0='d53465;
#10 word0='d53502;
#10 word0='d53539;
#10 word0='d53576;
#10 word0='d53613;
#10 word0='d53650;
#10 word0='d53687;
#10 word0='d53724;
#10 word0='d53761;
#10 word0='d53798;
#10 word0='d53835;
#10 word0='d53872;
#10 word0='d53909;
#10 word0='d53946;
#10 word0='d53983;
#10 word0='d54020;
#10 word0='d54057;
#10 word0='d54094;
#10 word0='d54131;
#10 word0='d54168;
#10 word0='d54205;
#10 word0='d54242;
#10 word0='d54279;
#10 word0='d54316;
#10 word0='d54353;
#10 word0='d54390;
#10 word0='d54427;
#10 word0='d54464;
#10 word0='d54501;
#10 word0='d54538;
#10 word0='d54575;
#10 word0='d54612;
#10 word0='d54649;
#10 word0='d54686;
#10 word0='d54723;
#10 word0='d54760;
#10 word0='d54797;
#10 word0='d54834;
#10 word0='d54871;
#10 word0='d54908;
#10 word0='d54945;
#10 word0='d54982;
#10 word0='d55019;
#10 word0='d55056;
#10 word0='d55093;
#10 word0='d55130;
#10 word0='d55167;
#10 word0='d55204;
#10 word0='d55241;
#10 word0='d55278;
#10 word0='d55315;
#10 word0='d55352;
#10 word0='d55389;
#10 word0='d55426;
#10 word0='d55463;
#10 word0='d55500;
#10 word0='d55537;
#10 word0='d55574;
#10 word0='d55611;
#10 word0='d55648;
#10 word0='d55685;
#10 word0='d55722;
#10 word0='d55759;
#10 word0='d55796;
#10 word0='d55833;
#10 word0='d55870;
#10 word0='d55907;
#10 word0='d55944;
#10 word0='d55981;
#10 word0='d56018;
#10 word0='d56055;
#10 word0='d56092;
#10 word0='d56129;
#10 word0='d56166;
#10 word0='d56203;
#10 word0='d56240;
#10 word0='d56277;
#10 word0='d56314;
#10 word0='d56351;
#10 word0='d56388;
#10 word0='d56425;
#10 word0='d56462;
#10 word0='d56499;
#10 word0='d56536;
#10 word0='d56573;
#10 word0='d56610;
#10 word0='d56647;
#10 word0='d56684;
#10 word0='d56721;
#10 word0='d56758;
#10 word0='d56795;
#10 word0='d56832;
#10 word0='d56869;
#10 word0='d56906;
#10 word0='d56943;
#10 word0='d56980;
#10 word0='d57017;
#10 word0='d57054;
#10 word0='d57091;
#10 word0='d57128;
#10 word0='d57165;
#10 word0='d57202;
#10 word0='d57239;
#10 word0='d57276;
#10 word0='d57313;
#10 word0='d57350;
#10 word0='d57387;
#10 word0='d57424;
#10 word0='d57461;
#10 word0='d57498;
#10 word0='d57535;
#10 word0='d57572;
#10 word0='d57609;
#10 word0='d57646;
#10 word0='d57683;
#10 word0='d57720;
#10 word0='d57757;
#10 word0='d57794;
#10 word0='d57831;
#10 word0='d57868;
#10 word0='d57905;
#10 word0='d57942;
#10 word0='d57979;
#10 word0='d58016;
#10 word0='d58053;
#10 word0='d58090;
#10 word0='d58127;
#10 word0='d58164;
#10 word0='d58201;
#10 word0='d58238;
#10 word0='d58275;
#10 word0='d58312;
#10 word0='d58349;
#10 word0='d58386;
#10 word0='d58423;
#10 word0='d58460;
#10 word0='d58497;
#10 word0='d58534;
#10 word0='d58571;
#10 word0='d58608;
#10 word0='d58645;
#10 word0='d58682;
#10 word0='d58719;
#10 word0='d58756;
#10 word0='d58793;
#10 word0='d58830;
#10 word0='d58867;
#10 word0='d58904;
#10 word0='d58941;
#10 word0='d58978;
#10 word0='d59015;
#10 word0='d59052;
#10 word0='d59089;
#10 word0='d59126;
#10 word0='d59163;
#10 word0='d59200;
#10 word0='d59237;
#10 word0='d59274;
#10 word0='d59311;
#10 word0='d59348;
#10 word0='d59385;
#10 word0='d59422;
#10 word0='d59459;
#10 word0='d59496;
#10 word0='d59533;
#10 word0='d59570;
#10 word0='d59607;
#10 word0='d59644;
#10 word0='d59681;
#10 word0='d59718;
#10 word0='d59755;
#10 word0='d59792;
#10 word0='d59829;
#10 word0='d59866;
#10 word0='d59903;
#10 word0='d59940;
#10 word0='d59977;
#10 word0='d60014;
#10 word0='d60051;
#10 word0='d60088;
#10 word0='d60125;
#10 word0='d60162;
#10 word0='d60199;
#10 word0='d60236;
#10 word0='d60273;
#10 word0='d60310;
#10 word0='d60347;
#10 word0='d60384;
#10 word0='d60421;
#10 word0='d60458;
#10 word0='d60495;
#10 word0='d60532;
#10 word0='d60569;
#10 word0='d60606;
#10 word0='d60643;
#10 word0='d60680;
#10 word0='d60717;
#10 word0='d60754;
#10 word0='d60791;
#10 word0='d60828;
#10 word0='d60865;
#10 word0='d60902;
#10 word0='d60939;
#10 word0='d60976;
#10 word0='d61013;
#10 word0='d61050;
#10 word0='d61087;
#10 word0='d61124;
#10 word0='d61161;
#10 word0='d61198;
#10 word0='d61235;
#10 word0='d61272;
#10 word0='d61309;
#10 word0='d61346;
#10 word0='d61383;
#10 word0='d61420;
#10 word0='d61457;
#10 word0='d61494;
#10 word0='d61531;
#10 word0='d61568;
#10 word0='d61605;
#10 word0='d61642;
#10 word0='d61679;
#10 word0='d61716;
#10 word0='d61753;
#10 word0='d61790;
#10 word0='d61827;
#10 word0='d61864;
#10 word0='d61901;
#10 word0='d61938;
#10 word0='d61975;
#10 word0='d62012;
#10 word0='d62049;
#10 word0='d62086;
#10 word0='d62123;
#10 word0='d62160;
#10 word0='d62197;
#10 word0='d62234;
#10 word0='d62271;
#10 word0='d62308;
#10 word0='d62345;
#10 word0='d62382;
#10 word0='d62419;
#10 word0='d62456;
#10 word0='d62493;
#10 word0='d62530;
#10 word0='d62567;
#10 word0='d62604;
#10 word0='d62641;
#10 word0='d62678;
#10 word0='d62715;
#10 word0='d62752;
#10 word0='d62789;
#10 word0='d62826;
#10 word0='d62863;
#10 word0='d62900;
#10 word0='d62937;
#10 word0='d62974;
#10 word0='d63011;
#10 word0='d63048;
#10 word0='d63085;
#10 word0='d63122;
#10 word0='d63159;
#10 word0='d63196;
#10 word0='d63233;
#10 word0='d63270;
#10 word0='d63307;
#10 word0='d63344;
#10 word0='d63381;
#10 word0='d63418;
#10 word0='d63455;
#10 word0='d63492;
#10 word0='d63529;
#10 word0='d63566;
#10 word0='d63603;
#10 word0='d63640;
#10 word0='d63677;
#10 word0='d63714;
#10 word0='d63751;
#10 word0='d63788;
#10 word0='d63825;
#10 word0='d63862;
#10 word0='d63899;
#10 word0='d63936;
#10 word0='d63973;
#10 word0='d64010;
#10 word0='d64047;
#10 word0='d64084;
#10 word0='d64121;
#10 word0='d64158;
#10 word0='d64195;
#10 word0='d64232;
#10 word0='d64269;
#10 word0='d64306;
#10 word0='d64343;
#10 word0='d64380;
#10 word0='d64417;
#10 word0='d64454;
#10 word0='d64491;
#10 word0='d64528;
#10 word0='d64565;
#10 word0='d64602;
#10 word0='d64639;
#10 word0='d64676;
#10 word0='d64713;
#10 word0='d64750;
#10 word0='d64787;
#10 word0='d64824;
#10 word0='d64861;
#10 word0='d64898;
#10 word0='d64935;
#10 word0='d64972;
#10 word0='d65009;
#10 word0='d65046;
#10 word0='d65083;
#10 word0='d65120;
#10 word0='d65157;
#10 word0='d65194;
#10 word0='d65231;
#10 word0='d65268;
#10 word0='d65305;
#10 word0='d65342;
#10 word0='d65379;
#10 word0='d65416;
#10 word0='d65453;
#10 word0='d65490;
#10 word0='d65527;
#10 word0='d65564;
#10 word0='d65601;
#10 word0='d65638;
#10 word0='d65675;
#10 word0='d65712;
#10 word0='d65749;
#10 word0='d65786;
#10 word0='d65823;
#10 word0='d65860;
#10 word0='d65897;
#10 word0='d65934;
#10 word0='d65971;
#10 word0='d66008;
#10 word0='d66045;
#10 word0='d66082;
#10 word0='d66119;
#10 word0='d66156;
#10 word0='d66193;
#10 word0='d66230;
#10 word0='d66267;
#10 word0='d66304;
#10 word0='d66341;
#10 word0='d66378;
#10 word0='d66415;
#10 word0='d66452;
#10 word0='d66489;
#10 word0='d66526;
#10 word0='d66563;
#10 word0='d66600;
#10 word0='d66637;
#10 word0='d66674;
#10 word0='d66711;
#10 word0='d66748;
#10 word0='d66785;
#10 word0='d66822;
#10 word0='d66859;
#10 word0='d66896;
#10 word0='d66933;
#10 word0='d66970;
#10 word0='d67007;
#10 word0='d67044;
#10 word0='d67081;
#10 word0='d67118;
#10 word0='d67155;
#10 word0='d67192;
#10 word0='d67229;
#10 word0='d67266;
#10 word0='d67303;
#10 word0='d67340;
#10 word0='d67377;
#10 word0='d67414;
#10 word0='d67451;
#10 word0='d67488;
#10 word0='d67525;
#10 word0='d67562;
#10 word0='d67599;
#10 word0='d67636;
#10 word0='d67673;
#10 word0='d67710;
#10 word0='d67747;
#10 word0='d67784;
#10 word0='d67821;
#10 word0='d67858;
#10 word0='d67895;
#10 word0='d67932;
#10 word0='d67969;
#10 word0='d68006;
#10 word0='d68043;
#10 word0='d68080;
#10 word0='d68117;
#10 word0='d68154;
#10 word0='d68191;
#10 word0='d68228;
#10 word0='d68265;
#10 word0='d68302;
#10 word0='d68339;
#10 word0='d68376;
#10 word0='d68413;
#10 word0='d68450;
#10 word0='d68487;
#10 word0='d68524;
#10 word0='d68561;
#10 word0='d68598;
#10 word0='d68635;
#10 word0='d68672;
#10 word0='d68709;
#10 word0='d68746;
#10 word0='d68783;
#10 word0='d68820;
#10 word0='d68857;
#10 word0='d68894;
#10 word0='d68931;
#10 word0='d68968;
#10 word0='d69005;
#10 word0='d69042;
#10 word0='d69079;
#10 word0='d69116;
#10 word0='d69153;
#10 word0='d69190;
#10 word0='d69227;
#10 word0='d69264;
#10 word0='d69301;
#10 word0='d69338;
#10 word0='d69375;
#10 word0='d69412;
#10 word0='d69449;
#10 word0='d69486;
#10 word0='d69523;
#10 word0='d69560;
#10 word0='d69597;
#10 word0='d69634;
#10 word0='d69671;
#10 word0='d69708;
#10 word0='d69745;
#10 word0='d69782;
#10 word0='d69819;
#10 word0='d69856;
#10 word0='d69893;
#10 word0='d69930;
#10 word0='d69967;
#10 word0='d70004;
#10 word0='d70041;
#10 word0='d70078;
#10 word0='d70115;
#10 word0='d70152;
#10 word0='d70189;
#10 word0='d70226;
#10 word0='d70263;
#10 word0='d70300;
#10 word0='d70337;
#10 word0='d70374;
#10 word0='d70411;
#10 word0='d70448;
#10 word0='d70485;
#10 word0='d70522;
#10 word0='d70559;
#10 word0='d70596;
#10 word0='d70633;
#10 word0='d70670;
#10 word0='d70707;
#10 word0='d70744;
#10 word0='d70781;
#10 word0='d70818;
#10 word0='d70855;
#10 word0='d70892;
#10 word0='d70929;
#10 word0='d70966;
#10 word0='d71003;
#10 word0='d71040;
#10 word0='d71077;
#10 word0='d71114;
#10 word0='d71151;
#10 word0='d71188;
#10 word0='d71225;
#10 word0='d71262;
#10 word0='d71299;
#10 word0='d71336;
#10 word0='d71373;
#10 word0='d71410;
#10 word0='d71447;
#10 word0='d71484;
#10 word0='d71521;
#10 word0='d71558;
#10 word0='d71595;
#10 word0='d71632;
#10 word0='d71669;
#10 word0='d71706;
#10 word0='d71743;
#10 word0='d71780;
#10 word0='d71817;
#10 word0='d71854;
#10 word0='d71891;
#10 word0='d71928;
#10 word0='d71965;
#10 word0='d72002;
#10 word0='d72039;
#10 word0='d72076;
#10 word0='d72113;
#10 word0='d72150;
#10 word0='d72187;
#10 word0='d72224;
#10 word0='d72261;
#10 word0='d72298;
#10 word0='d72335;
#10 word0='d72372;
#10 word0='d72409;
#10 word0='d72446;
#10 word0='d72483;
#10 word0='d72520;
#10 word0='d72557;
#10 word0='d72594;
#10 word0='d72631;
#10 word0='d72668;
#10 word0='d72705;
#10 word0='d72742;
#10 word0='d72779;
#10 word0='d72816;
#10 word0='d72853;
#10 word0='d72890;
#10 word0='d72927;
#10 word0='d72964;
#10 word0='d73001;
#10 word0='d73038;
#10 word0='d73075;
#10 word0='d73112;
#10 word0='d73149;
#10 word0='d73186;
#10 word0='d73223;
#10 word0='d73260;
#10 word0='d73297;
#10 word0='d73334;
#10 word0='d73371;
#10 word0='d73408;
#10 word0='d73445;
#10 word0='d73482;
#10 word0='d73519;
#10 word0='d73556;
#10 word0='d73593;
#10 word0='d73630;
#10 word0='d73667;
#10 word0='d73704;
#10 word0='d73741;
#10 word0='d73778;
#10 word0='d73815;
#10 word0='d73852;
#10 word0='d73889;
#10 word0='d73926;
#10 word0='d73963;
#10 word0='d74000;
#10 word0='d74037;
#10 word0='d74074;
#10 word0='d74111;
#10 word0='d74148;
#10 word0='d74185;
#10 word0='d74222;
#10 word0='d74259;
#10 word0='d74296;
#10 word0='d74333;
#10 word0='d74370;
#10 word0='d74407;
#10 word0='d74444;
#10 word0='d74481;
#10 word0='d74518;
#10 word0='d74555;
#10 word0='d74592;
#10 word0='d74629;
#10 word0='d74666;
#10 word0='d74703;
#10 word0='d74740;
#10 word0='d74777;
#10 word0='d74814;
#10 word0='d74851;
#10 word0='d74888;
#10 word0='d74925;
#10 word0='d74962;
#10 word0='d74999;
#10 word0='d75036;
#10 word0='d75073;
#10 word0='d75110;
#10 word0='d75147;
#10 word0='d75184;
#10 word0='d75221;
#10 word0='d75258;
#10 word0='d75295;
#10 word0='d75332;
#10 word0='d75369;
#10 word0='d75406;
#10 word0='d75443;
#10 word0='d75480;
#10 word0='d75517;
#10 word0='d75554;
#10 word0='d75591;
#10 word0='d75628;
#10 word0='d75665;
#10 word0='d75702;
#10 word0='d75739;
#10 word0='d75776;
#10 word0='d75813;
#10 word0='d75850;
#10 word0='d75887;
#10 word0='d75924;
#10 word0='d75961;
#10 word0='d75998;
#10 word0='d76035;
#10 word0='d76072;
#10 word0='d76109;
#10 word0='d76146;
#10 word0='d76183;
#10 word0='d76220;
#10 word0='d76257;
#10 word0='d76294;
#10 word0='d76331;
#10 word0='d76368;
#10 word0='d76405;
#10 word0='d76442;
#10 word0='d76479;
#10 word0='d76516;
#10 word0='d76553;
#10 word0='d76590;
#10 word0='d76627;
#10 word0='d76664;
#10 word0='d76701;
#10 word0='d76738;
#10 word0='d76775;
#10 word0='d76812;
#10 word0='d76849;
#10 word0='d76886;
#10 word0='d76923;
#10 word0='d76960;
#10 word0='d76997;
#10 word0='d77034;
#10 word0='d77071;
#10 word0='d77108;
#10 word0='d77145;
#10 word0='d77182;
#10 word0='d77219;
#10 word0='d77256;
#10 word0='d77293;
#10 word0='d77330;
#10 word0='d77367;
#10 word0='d77404;
#10 word0='d77441;
#10 word0='d77478;
#10 word0='d77515;
#10 word0='d77552;
#10 word0='d77589;
#10 word0='d77626;
#10 word0='d77663;
#10 word0='d77700;
#10 word0='d77737;
#10 word0='d77774;
#10 word0='d77811;
#10 word0='d77848;
#10 word0='d77885;
#10 word0='d77922;
#10 word0='d77959;
#10 word0='d77996;
#10 word0='d78033;
#10 word0='d78070;
#10 word0='d78107;
#10 word0='d78144;
#10 word0='d78181;
#10 word0='d78218;
#10 word0='d78255;
#10 word0='d78292;
#10 word0='d78329;
#10 word0='d78366;
#10 word0='d78403;
#10 word0='d78440;
#10 word0='d78477;
#10 word0='d78514;
#10 word0='d78551;
#10 word0='d78588;
#10 word0='d78625;
#10 word0='d78662;
#10 word0='d78699;
#10 word0='d78736;
#10 word0='d78773;
#10 word0='d78810;
#10 word0='d78847;
#10 word0='d78884;
#10 word0='d78921;
#10 word0='d78958;
#10 word0='d78995;
#10 word0='d79032;
#10 word0='d79069;
#10 word0='d79106;
#10 word0='d79143;
#10 word0='d79180;
#10 word0='d79217;
#10 word0='d79254;
#10 word0='d79291;
#10 word0='d79328;
#10 word0='d79365;
#10 word0='d79402;
#10 word0='d79439;
#10 word0='d79476;
#10 word0='d79513;
#10 word0='d79550;
#10 word0='d79587;
#10 word0='d79624;
#10 word0='d79661;
#10 word0='d79698;
#10 word0='d79735;
#10 word0='d79772;
#10 word0='d79809;
#10 word0='d79846;
#10 word0='d79883;
#10 word0='d79920;
#10 word0='d79957;
#10 word0='d79994;
#10 word0='d80031;
#10 word0='d80068;
#10 word0='d80105;
#10 word0='d80142;
#10 word0='d80179;
#10 word0='d80216;
#10 word0='d80253;
#10 word0='d80290;
#10 word0='d80327;
#10 word0='d80364;
#10 word0='d80401;
#10 word0='d80438;
#10 word0='d80475;
#10 word0='d80512;
#10 word0='d80549;
#10 word0='d80586;
#10 word0='d80623;
#10 word0='d80660;
#10 word0='d80697;
#10 word0='d80734;
#10 word0='d80771;
#10 word0='d80808;
#10 word0='d80845;
#10 word0='d80882;
#10 word0='d80919;
#10 word0='d80956;
#10 word0='d80993;
#10 word0='d81030;
#10 word0='d81067;
#10 word0='d81104;
#10 word0='d81141;
#10 word0='d81178;
#10 word0='d81215;
#10 word0='d81252;
#10 word0='d81289;
#10 word0='d81326;
#10 word0='d81363;
#10 word0='d81400;
#10 word0='d81437;
#10 word0='d81474;
#10 word0='d81511;
#10 word0='d81548;
#10 word0='d81585;
#10 word0='d81622;
#10 word0='d81659;
#10 word0='d81696;
#10 word0='d81733;
#10 word0='d81770;
#10 word0='d81807;
#10 word0='d81844;
#10 word0='d81881;
#10 word0='d81918;
#10 word0='d81955;
#10 word0='d81992;
#10 word0='d82029;
#10 word0='d82066;
#10 word0='d82103;
#10 word0='d82140;
#10 word0='d82177;
#10 word0='d82214;
#10 word0='d82251;
#10 word0='d82288;
#10 word0='d82325;
#10 word0='d82362;
#10 word0='d82399;
#10 word0='d82436;
#10 word0='d82473;
#10 word0='d82510;
#10 word0='d82547;
#10 word0='d82584;
#10 word0='d82621;
#10 word0='d82658;
#10 word0='d82695;
#10 word0='d82732;
#10 word0='d82769;
#10 word0='d82806;
#10 word0='d82843;
#10 word0='d82880;
#10 word0='d82917;
#10 word0='d82954;
#10 word0='d82991;
#10 word0='d83028;
#10 word0='d83065;
#10 word0='d83102;
#10 word0='d83139;
#10 word0='d83176;
#10 word0='d83213;
#10 word0='d83250;
#10 word0='d83287;
#10 word0='d83324;
#10 word0='d83361;
#10 word0='d83398;
#10 word0='d83435;
#10 word0='d83472;
#10 word0='d83509;
#10 word0='d83546;
#10 word0='d83583;
#10 word0='d83620;
#10 word0='d83657;
#10 word0='d83694;
#10 word0='d83731;
#10 word0='d83768;
#10 word0='d83805;
#10 word0='d83842;
#10 word0='d83879;
#10 word0='d83916;
#10 word0='d83953;
#10 word0='d83990;
#10 word0='d84027;
#10 word0='d84064;
#10 word0='d84101;
#10 word0='d84138;
#10 word0='d84175;
#10 word0='d84212;
#10 word0='d84249;
#10 word0='d84286;
#10 word0='d84323;
#10 word0='d84360;
#10 word0='d84397;
#10 word0='d84434;
#10 word0='d84471;
#10 word0='d84508;
#10 word0='d84545;
#10 word0='d84582;
#10 word0='d84619;
#10 word0='d84656;
#10 word0='d84693;
#10 word0='d84730;
#10 word0='d84767;
#10 word0='d84804;
#10 word0='d84841;
#10 word0='d84878;
#10 word0='d84915;
#10 word0='d84952;
#10 word0='d84989;
#10 word0='d85026;
#10 word0='d85063;
#10 word0='d85100;
#10 word0='d85137;
#10 word0='d85174;
#10 word0='d85211;
#10 word0='d85248;
#10 word0='d85285;
#10 word0='d85322;
#10 word0='d85359;
#10 word0='d85396;
#10 word0='d85433;
#10 word0='d85470;
#10 word0='d85507;
#10 word0='d85544;
#10 word0='d85581;
#10 word0='d85618;
#10 word0='d85655;
#10 word0='d85692;
#10 word0='d85729;
#10 word0='d85766;
#10 word0='d85803;
#10 word0='d85840;
#10 word0='d85877;
#10 word0='d85914;
#10 word0='d85951;
#10 word0='d85988;
#10 word0='d86025;
#10 word0='d86062;
#10 word0='d86099;
#10 word0='d86136;
#10 word0='d86173;
#10 word0='d86210;
#10 word0='d86247;
#10 word0='d86284;
#10 word0='d86321;
#10 word0='d86358;
#10 word0='d86395;
#10 word0='d86432;
#10 word0='d86469;
#10 word0='d86506;
#10 word0='d86543;
#10 word0='d86580;
#10 word0='d86617;
#10 word0='d86654;
#10 word0='d86691;
#10 word0='d86728;
#10 word0='d86765;
#10 word0='d86802;
#10 word0='d86839;
#10 word0='d86876;
#10 word0='d86913;
#10 word0='d86950;
#10 word0='d86987;
#10 word0='d87024;
#10 word0='d87061;
#10 word0='d87098;
#10 word0='d87135;
#10 word0='d87172;
#10 word0='d87209;
#10 word0='d87246;
#10 word0='d87283;
#10 word0='d87320;
#10 word0='d87357;
#10 word0='d87394;
#10 word0='d87431;
#10 word0='d87468;
#10 word0='d87505;
#10 word0='d87542;
#10 word0='d87579;
#10 word0='d87616;
#10 word0='d87653;
#10 word0='d87690;
#10 word0='d87727;
#10 word0='d87764;
#10 word0='d87801;
#10 word0='d87838;
#10 word0='d87875;
#10 word0='d87912;
#10 word0='d87949;
#10 word0='d87986;
#10 word0='d88023;
#10 word0='d88060;
#10 word0='d88097;
#10 word0='d88134;
#10 word0='d88171;
#10 word0='d88208;
#10 word0='d88245;
#10 word0='d88282;
#10 word0='d88319;
#10 word0='d88356;
#10 word0='d88393;
#10 word0='d88430;
#10 word0='d88467;
#10 word0='d88504;
#10 word0='d88541;
#10 word0='d88578;
#10 word0='d88615;
#10 word0='d88652;
#10 word0='d88689;
#10 word0='d88726;
#10 word0='d88763;
#10 word0='d88800;
#10 word0='d88837;
#10 word0='d88874;
#10 word0='d88911;
#10 word0='d88948;
#10 word0='d88985;
#10 word0='d89022;
#10 word0='d89059;
#10 word0='d89096;
#10 word0='d89133;
#10 word0='d89170;
#10 word0='d89207;
#10 word0='d89244;
#10 word0='d89281;
#10 word0='d89318;
#10 word0='d89355;
#10 word0='d89392;
#10 word0='d89429;
#10 word0='d89466;
#10 word0='d89503;
#10 word0='d89540;
#10 word0='d89577;
#10 word0='d89614;
#10 word0='d89651;
#10 word0='d89688;
#10 word0='d89725;
#10 word0='d89762;
#10 word0='d89799;
#10 word0='d89836;
#10 word0='d89873;
#10 word0='d89910;
#10 word0='d89947;
#10 word0='d89984;
#10 word0='d90021;
#10 word0='d90058;
#10 word0='d90095;
#10 word0='d90132;
#10 word0='d90169;
#10 word0='d90206;
#10 word0='d90243;
#10 word0='d90280;
#10 word0='d90317;
#10 word0='d90354;
#10 word0='d90391;
#10 word0='d90428;
#10 word0='d90465;
#10 word0='d90502;
#10 word0='d90539;
#10 word0='d90576;
#10 word0='d90613;
#10 word0='d90650;
#10 word0='d90687;
#10 word0='d90724;
#10 word0='d90761;
#10 word0='d90798;
#10 word0='d90835;
#10 word0='d90872;
#10 word0='d90909;
#10 word0='d90946;
#10 word0='d90983;
#10 word0='d91020;
#10 word0='d91057;
#10 word0='d91094;
#10 word0='d91131;
#10 word0='d91168;
#10 word0='d91205;
#10 word0='d91242;
#10 word0='d91279;
#10 word0='d91316;
#10 word0='d91353;
#10 word0='d91390;
#10 word0='d91427;
#10 word0='d91464;
#10 word0='d91501;
#10 word0='d91538;
#10 word0='d91575;
#10 word0='d91612;
#10 word0='d91649;
#10 word0='d91686;
#10 word0='d91723;
#10 word0='d91760;
#10 word0='d91797;
#10 word0='d91834;
#10 word0='d91871;
#10 word0='d91908;
#10 word0='d91945;
#10 word0='d91982;
#10 word0='d92019;
#10 word0='d92056;
#10 word0='d92093;
#10 word0='d92130;
#10 word0='d92167;
#10 word0='d92204;
#10 word0='d92241;
#10 word0='d92278;
#10 word0='d92315;
#10 word0='d92352;
#10 word0='d92389;
#10 word0='d92426;
#10 word0='d92463;
#10 word0='d92500;
#10 word0='d92537;
#10 word0='d92574;
#10 word0='d92611;
#10 word0='d92648;
#10 word0='d92685;
#10 word0='d92722;
#10 word0='d92759;
#10 word0='d92796;
#10 word0='d92833;
#10 word0='d92870;
#10 word0='d92907;
#10 word0='d92944;
#10 word0='d92981;
#10 word0='d93018;
#10 word0='d93055;
#10 word0='d93092;
#10 word0='d93129;
#10 word0='d93166;
#10 word0='d93203;
#10 word0='d93240;
#10 word0='d93277;
#10 word0='d93314;
#10 word0='d93351;
#10 word0='d93388;
#10 word0='d93425;
#10 word0='d93462;
#10 word0='d93499;
#10 word0='d93536;
#10 word0='d93573;
#10 word0='d93610;
#10 word0='d93647;
#10 word0='d93684;
#10 word0='d93721;
#10 word0='d93758;
#10 word0='d93795;
#10 word0='d93832;
#10 word0='d93869;
#10 word0='d93906;
#10 word0='d93943;
#10 word0='d93980;
#10 word0='d94017;
#10 word0='d94054;
#10 word0='d94091;
#10 word0='d94128;
#10 word0='d94165;
#10 word0='d94202;
#10 word0='d94239;
#10 word0='d94276;
#10 word0='d94313;
#10 word0='d94350;
#10 word0='d94387;
#10 word0='d94424;
#10 word0='d94461;
#10 word0='d94498;
#10 word0='d94535;
#10 word0='d94572;
#10 word0='d94609;
#10 word0='d94646;
#10 word0='d94683;
#10 word0='d94720;
#10 word0='d94757;
#10 word0='d94794;
#10 word0='d94831;
#10 word0='d94868;
#10 word0='d94905;
#10 word0='d94942;
#10 word0='d94979;
#10 word0='d95016;
#10 word0='d95053;
#10 word0='d95090;
#10 word0='d95127;
#10 word0='d95164;
#10 word0='d95201;
#10 word0='d95238;
#10 word0='d95275;
#10 word0='d95312;
#10 word0='d95349;
#10 word0='d95386;
#10 word0='d95423;
#10 word0='d95460;
#10 word0='d95497;
#10 word0='d95534;
#10 word0='d95571;
#10 word0='d95608;
#10 word0='d95645;
#10 word0='d95682;
#10 word0='d95719;
#10 word0='d95756;
#10 word0='d95793;
#10 word0='d95830;
#10 word0='d95867;
#10 word0='d95904;
#10 word0='d95941;
#10 word0='d95978;
#10 word0='d96015;
#10 word0='d96052;
#10 word0='d96089;
#10 word0='d96126;
#10 word0='d96163;
#10 word0='d96200;
#10 word0='d96237;
#10 word0='d96274;
#10 word0='d96311;
#10 word0='d96348;
#10 word0='d96385;
#10 word0='d96422;
#10 word0='d96459;
#10 word0='d96496;
#10 word0='d96533;
#10 word0='d96570;
#10 word0='d96607;
#10 word0='d96644;
#10 word0='d96681;
#10 word0='d96718;
#10 word0='d96755;
#10 word0='d96792;
#10 word0='d96829;
#10 word0='d96866;
#10 word0='d96903;
#10 word0='d96940;
#10 word0='d96977;
#10 word0='d97014;
#10 word0='d97051;
#10 word0='d97088;
#10 word0='d97125;
#10 word0='d97162;
#10 word0='d97199;
#10 word0='d97236;
#10 word0='d97273;
#10 word0='d97310;
#10 word0='d97347;
#10 word0='d97384;
#10 word0='d97421;
#10 word0='d97458;
#10 word0='d97495;
#10 word0='d97532;
#10 word0='d97569;
#10 word0='d97606;
#10 word0='d97643;
#10 word0='d97680;
#10 word0='d97717;
#10 word0='d97754;
#10 word0='d97791;
#10 word0='d97828;
#10 word0='d97865;
#10 word0='d97902;
#10 word0='d97939;
#10 word0='d97976;
#10 word0='d98013;
#10 word0='d98050;
#10 word0='d98087;
#10 word0='d98124;
#10 word0='d98161;
#10 word0='d98198;
#10 word0='d98235;
#10 word0='d98272;
#10 word0='d98309;
#10 word0='d98346;
#10 word0='d98383;
#10 word0='d98420;
#10 word0='d98457;
#10 word0='d98494;
#10 word0='d98531;
#10 word0='d98568;
#10 word0='d98605;
#10 word0='d98642;
#10 word0='d98679;
#10 word0='d98716;
#10 word0='d98753;
#10 word0='d98790;
#10 word0='d98827;
#10 word0='d98864;
#10 word0='d98901;
#10 word0='d98938;
#10 word0='d98975;
#10 word0='d99012;
#10 word0='d99049;
#10 word0='d99086;
#10 word0='d99123;
#10 word0='d99160;
#10 word0='d99197;
#10 word0='d99234;
#10 word0='d99271;
#10 word0='d99308;
#10 word0='d99345;
#10 word0='d99382;
#10 word0='d99419;
#10 word0='d99456;
#10 word0='d99493;
#10 word0='d99530;
#10 word0='d99567;
#10 word0='d99604;
#10 word0='d99641;
#10 word0='d99678;
#10 word0='d99715;
#10 word0='d99752;
#10 word0='d99789;
#10 word0='d99826;
#10 word0='d99863;
#10 word0='d99900;
#10 word0='d99937;
#10 word0='d99974;
#10 word0='d100011;
#10 word0='d100048;
#10 word0='d100085;
#10 word0='d100122;
#10 word0='d100159;
#10 word0='d100196;
#10 word0='d100233;
#10 word0='d100270;
#10 word0='d100307;
#10 word0='d100344;
#10 word0='d100381;
#10 word0='d100418;
#10 word0='d100455;
#10 word0='d100492;
#10 word0='d100529;
#10 word0='d100566;
#10 word0='d100603;
#10 word0='d100640;
#10 word0='d100677;
#10 word0='d100714;
#10 word0='d100751;
#10 word0='d100788;
#10 word0='d100825;
#10 word0='d100862;
#10 word0='d100899;
#10 word0='d100936;
#10 word0='d100973;
#10 word0='d101010;
#10 word0='d101047;
#10 word0='d101084;
#10 word0='d101121;
#10 word0='d101158;
#10 word0='d101195;
#10 word0='d101232;
#10 word0='d101269;
#10 word0='d101306;
#10 word0='d101343;
#10 word0='d101380;
#10 word0='d101417;
#10 word0='d101454;
#10 word0='d101491;
#10 word0='d101528;
#10 word0='d101565;
#10 word0='d101602;
#10 word0='d101639;
#10 word0='d101676;
#10 word0='d101713;
#10 word0='d101750;
#10 word0='d101787;
#10 word0='d101824;
#10 word0='d101861;
#10 word0='d101898;
#10 word0='d101935;
#10 word0='d101972;
#10 word0='d102009;
#10 word0='d102046;
#10 word0='d102083;
#10 word0='d102120;
#10 word0='d102157;
#10 word0='d102194;
#10 word0='d102231;
#10 word0='d102268;
#10 word0='d102305;
#10 word0='d102342;
#10 word0='d102379;
#10 word0='d102416;
#10 word0='d102453;
#10 word0='d102490;
#10 word0='d102527;
#10 word0='d102564;
#10 word0='d102601;
#10 word0='d102638;
#10 word0='d102675;
#10 word0='d102712;
#10 word0='d102749;
#10 word0='d102786;
#10 word0='d102823;
#10 word0='d102860;
#10 word0='d102897;
#10 word0='d102934;
#10 word0='d102971;
#10 word0='d103008;
#10 word0='d103045;
#10 word0='d103082;
#10 word0='d103119;
#10 word0='d103156;
#10 word0='d103193;
#10 word0='d103230;
#10 word0='d103267;
#10 word0='d103304;
#10 word0='d103341;
#10 word0='d103378;
#10 word0='d103415;
#10 word0='d103452;
#10 word0='d103489;
#10 word0='d103526;
#10 word0='d103563;
#10 word0='d103600;
#10 word0='d103637;
#10 word0='d103674;
#10 word0='d103711;
#10 word0='d103748;
#10 word0='d103785;
#10 word0='d103822;
#10 word0='d103859;
#10 word0='d103896;
#10 word0='d103933;
#10 word0='d103970;
#10 word0='d104007;
#10 word0='d104044;
#10 word0='d104081;
#10 word0='d104118;
#10 word0='d104155;
#10 word0='d104192;
#10 word0='d104229;
#10 word0='d104266;
#10 word0='d104303;
#10 word0='d104340;
#10 word0='d104377;
#10 word0='d104414;
#10 word0='d104451;
#10 word0='d104488;
#10 word0='d104525;
#10 word0='d104562;
#10 word0='d104599;
#10 word0='d104636;
#10 word0='d104673;
#10 word0='d104710;
#10 word0='d104747;
#10 word0='d104784;
#10 word0='d104821;
#10 word0='d104858;
#10 word0='d104895;
#10 word0='d104932;
#10 word0='d104969;
#10 word0='d105006;
#10 word0='d105043;
#10 word0='d105080;
#10 word0='d105117;
#10 word0='d105154;
#10 word0='d105191;
#10 word0='d105228;
#10 word0='d105265;
#10 word0='d105302;
#10 word0='d105339;
#10 word0='d105376;
#10 word0='d105413;
#10 word0='d105450;
#10 word0='d105487;
#10 word0='d105524;
#10 word0='d105561;
#10 word0='d105598;
#10 word0='d105635;
#10 word0='d105672;
#10 word0='d105709;
#10 word0='d105746;
#10 word0='d105783;
#10 word0='d105820;
#10 word0='d105857;
#10 word0='d105894;
#10 word0='d105931;
#10 word0='d105968;
#10 word0='d106005;
#10 word0='d106042;
#10 word0='d106079;
#10 word0='d106116;
#10 word0='d106153;
#10 word0='d106190;
#10 word0='d106227;
#10 word0='d106264;
#10 word0='d106301;
#10 word0='d106338;
#10 word0='d106375;
#10 word0='d106412;
#10 word0='d106449;
#10 word0='d106486;
#10 word0='d106523;
#10 word0='d106560;
#10 word0='d106597;
#10 word0='d106634;
#10 word0='d106671;
#10 word0='d106708;
#10 word0='d106745;
#10 word0='d106782;
#10 word0='d106819;
#10 word0='d106856;
#10 word0='d106893;
#10 word0='d106930;
#10 word0='d106967;
#10 word0='d107004;
#10 word0='d107041;
#10 word0='d107078;
#10 word0='d107115;
#10 word0='d107152;
#10 word0='d107189;
#10 word0='d107226;
#10 word0='d107263;
#10 word0='d107300;
#10 word0='d107337;
#10 word0='d107374;
#10 word0='d107411;
#10 word0='d107448;
#10 word0='d107485;
#10 word0='d107522;
#10 word0='d107559;
#10 word0='d107596;
#10 word0='d107633;
#10 word0='d107670;
#10 word0='d107707;
#10 word0='d107744;
#10 word0='d107781;
#10 word0='d107818;
#10 word0='d107855;
#10 word0='d107892;
#10 word0='d107929;
#10 word0='d107966;
#10 word0='d108003;
#10 word0='d108040;
#10 word0='d108077;
#10 word0='d108114;
#10 word0='d108151;
#10 word0='d108188;
#10 word0='d108225;
#10 word0='d108262;
#10 word0='d108299;
#10 word0='d108336;
#10 word0='d108373;
#10 word0='d108410;
#10 word0='d108447;
#10 word0='d108484;
#10 word0='d108521;
#10 word0='d108558;
#10 word0='d108595;
#10 word0='d108632;
#10 word0='d108669;
#10 word0='d108706;
#10 word0='d108743;
#10 word0='d108780;
#10 word0='d108817;
#10 word0='d108854;
#10 word0='d108891;
#10 word0='d108928;
#10 word0='d108965;
#10 word0='d109002;
#10 word0='d109039;
#10 word0='d109076;
#10 word0='d109113;
#10 word0='d109150;
#10 word0='d109187;
#10 word0='d109224;
#10 word0='d109261;
#10 word0='d109298;
#10 word0='d109335;
#10 word0='d109372;
#10 word0='d109409;
#10 word0='d109446;
#10 word0='d109483;
#10 word0='d109520;
#10 word0='d109557;
#10 word0='d109594;
#10 word0='d109631;
#10 word0='d109668;
#10 word0='d109705;
#10 word0='d109742;
#10 word0='d109779;
#10 word0='d109816;
#10 word0='d109853;
#10 word0='d109890;
#10 word0='d109927;
#10 word0='d109964;
#10 word0='d110001;
#10 word0='d110038;
#10 word0='d110075;
#10 word0='d110112;
#10 word0='d110149;
#10 word0='d110186;
#10 word0='d110223;
#10 word0='d110260;
#10 word0='d110297;
#10 word0='d110334;
#10 word0='d110371;
#10 word0='d110408;
#10 word0='d110445;
#10 word0='d110482;
#10 word0='d110519;
#10 word0='d110556;
#10 word0='d110593;
#10 word0='d110630;
#10 word0='d110667;
#10 word0='d110704;
#10 word0='d110741;
#10 word0='d110778;
#10 word0='d110815;
#10 word0='d110852;
#10 word0='d110889;
#10 word0='d110926;
#10 word0='d110963;
#10 word0='d111000;
#10 word0='d111037;
#10 word0='d111074;
#10 word0='d111111;
#10 word0='d111148;
#10 word0='d111185;
#10 word0='d111222;
#10 word0='d111259;
#10 word0='d111296;
#10 word0='d111333;
#10 word0='d111370;
#10 word0='d111407;
#10 word0='d111444;
#10 word0='d111481;
#10 word0='d111518;
#10 word0='d111555;
#10 word0='d111592;
#10 word0='d111629;
#10 word0='d111666;
#10 word0='d111703;
#10 word0='d111740;
#10 word0='d111777;
#10 word0='d111814;
#10 word0='d111851;
#10 word0='d111888;
#10 word0='d111925;
#10 word0='d111962;
#10 word0='d111999;
#10 word0='d112036;
#10 word0='d112073;
#10 word0='d112110;
#10 word0='d112147;
#10 word0='d112184;
#10 word0='d112221;
#10 word0='d112258;
#10 word0='d112295;
#10 word0='d112332;
#10 word0='d112369;
#10 word0='d112406;
#10 word0='d112443;
#10 word0='d112480;
#10 word0='d112517;
#10 word0='d112554;
#10 word0='d112591;
#10 word0='d112628;
#10 word0='d112665;
#10 word0='d112702;
#10 word0='d112739;
#10 word0='d112776;
#10 word0='d112813;
#10 word0='d112850;
#10 word0='d112887;
#10 word0='d112924;
#10 word0='d112961;
#10 word0='d112998;
#10 word0='d113035;
#10 word0='d113072;
#10 word0='d113109;
#10 word0='d113146;
#10 word0='d113183;
#10 word0='d113220;
#10 word0='d113257;
#10 word0='d113294;
#10 word0='d113331;
#10 word0='d113368;
#10 word0='d113405;
#10 word0='d113442;
#10 word0='d113479;
#10 word0='d113516;
#10 word0='d113553;
#10 word0='d113590;
#10 word0='d113627;
#10 word0='d113664;
#10 word0='d113701;
#10 word0='d113738;
#10 word0='d113775;
#10 word0='d113812;
#10 word0='d113849;
#10 word0='d113886;
#10 word0='d113923;
#10 word0='d113960;
#10 word0='d113997;
#10 word0='d114034;
#10 word0='d114071;
#10 word0='d114108;
#10 word0='d114145;
#10 word0='d114182;
#10 word0='d114219;
#10 word0='d114256;
#10 word0='d114293;
#10 word0='d114330;
#10 word0='d114367;
#10 word0='d114404;
#10 word0='d114441;
#10 word0='d114478;
#10 word0='d114515;
#10 word0='d114552;
#10 word0='d114589;
#10 word0='d114626;
#10 word0='d114663;
#10 word0='d114700;
#10 word0='d114737;
#10 word0='d114774;
#10 word0='d114811;
#10 word0='d114848;
#10 word0='d114885;
#10 word0='d114922;
#10 word0='d114959;
#10 word0='d114996;
#10 word0='d115033;
#10 word0='d115070;
#10 word0='d115107;
#10 word0='d115144;
#10 word0='d115181;
#10 word0='d115218;
#10 word0='d115255;
#10 word0='d115292;
#10 word0='d115329;
#10 word0='d115366;
#10 word0='d115403;
#10 word0='d115440;
#10 word0='d115477;
#10 word0='d115514;
#10 word0='d115551;
#10 word0='d115588;
#10 word0='d115625;
#10 word0='d115662;
#10 word0='d115699;
#10 word0='d115736;
#10 word0='d115773;
#10 word0='d115810;
#10 word0='d115847;
#10 word0='d115884;
#10 word0='d115921;
#10 word0='d115958;
#10 word0='d115995;
#10 word0='d116032;
#10 word0='d116069;
#10 word0='d116106;
#10 word0='d116143;
#10 word0='d116180;
#10 word0='d116217;
#10 word0='d116254;
#10 word0='d116291;
#10 word0='d116328;
#10 word0='d116365;
#10 word0='d116402;
#10 word0='d116439;
#10 word0='d116476;
#10 word0='d116513;
#10 word0='d116550;
#10 word0='d116587;
#10 word0='d116624;
#10 word0='d116661;
#10 word0='d116698;
#10 word0='d116735;
#10 word0='d116772;
#10 word0='d116809;
#10 word0='d116846;
#10 word0='d116883;
#10 word0='d116920;
#10 word0='d116957;
#10 word0='d116994;
#10 word0='d117031;
#10 word0='d117068;
#10 word0='d117105;
#10 word0='d117142;
#10 word0='d117179;
#10 word0='d117216;
#10 word0='d117253;
#10 word0='d117290;
#10 word0='d117327;
#10 word0='d117364;
#10 word0='d117401;
#10 word0='d117438;
#10 word0='d117475;
#10 word0='d117512;
#10 word0='d117549;
#10 word0='d117586;
#10 word0='d117623;
#10 word0='d117660;
#10 word0='d117697;
#10 word0='d117734;
#10 word0='d117771;
#10 word0='d117808;
#10 word0='d117845;
#10 word0='d117882;
#10 word0='d117919;
#10 word0='d117956;
#10 word0='d117993;
#10 word0='d118030;
#10 word0='d118067;
#10 word0='d118104;
#10 word0='d118141;
#10 word0='d118178;
#10 word0='d118215;
#10 word0='d118252;
#10 word0='d118289;
#10 word0='d118326;
#10 word0='d118363;
#10 word0='d118400;
#10 word0='d118437;
#10 word0='d118474;
#10 word0='d118511;
#10 word0='d118548;
#10 word0='d118585;
#10 word0='d118622;
#10 word0='d118659;
#10 word0='d118696;
#10 word0='d118733;
#10 word0='d118770;
#10 word0='d118807;
#10 word0='d118844;
#10 word0='d118881;
#10 word0='d118918;
#10 word0='d118955;
#10 word0='d118992;
#10 word0='d119029;
#10 word0='d119066;
#10 word0='d119103;
#10 word0='d119140;
#10 word0='d119177;
#10 word0='d119214;
#10 word0='d119251;
#10 word0='d119288;
#10 word0='d119325;
#10 word0='d119362;
#10 word0='d119399;
#10 word0='d119436;
#10 word0='d119473;
#10 word0='d119510;
#10 word0='d119547;
#10 word0='d119584;
#10 word0='d119621;
#10 word0='d119658;
#10 word0='d119695;
#10 word0='d119732;
#10 word0='d119769;
#10 word0='d119806;
#10 word0='d119843;
#10 word0='d119880;
#10 word0='d119917;
#10 word0='d119954;
#10 word0='d119991;
#10 word0='d120028;
#10 word0='d120065;
#10 word0='d120102;
#10 word0='d120139;
#10 word0='d120176;
#10 word0='d120213;
#10 word0='d120250;
#10 word0='d120287;
#10 word0='d120324;
#10 word0='d120361;
#10 word0='d120398;
#10 word0='d120435;
#10 word0='d120472;
#10 word0='d120509;
#10 word0='d120546;
#10 word0='d120583;
#10 word0='d120620;
#10 word0='d120657;
#10 word0='d120694;
#10 word0='d120731;
#10 word0='d120768;
#10 word0='d120805;
#10 word0='d120842;
#10 word0='d120879;
#10 word0='d120916;
#10 word0='d120953;
#10 word0='d120990;
#10 word0='d121027;
#10 word0='d121064;
#10 word0='d121101;
#10 word0='d121138;
#10 word0='d121175;
#10 word0='d121212;
#10 word0='d121249;
#10 word0='d121286;
#10 word0='d121323;
#10 word0='d121360;
#10 word0='d121397;
#10 word0='d121434;
#10 word0='d121471;
#10 word0='d121508;
#10 word0='d121545;
#10 word0='d121582;
#10 word0='d121619;
#10 word0='d121656;
#10 word0='d121693;
#10 word0='d121730;
#10 word0='d121767;
#10 word0='d121804;
#10 word0='d121841;
#10 word0='d121878;
#10 word0='d121915;
#10 word0='d121952;
#10 word0='d121989;
#10 word0='d122026;
#10 word0='d122063;
#10 word0='d122100;
#10 word0='d122137;
#10 word0='d122174;
#10 word0='d122211;
#10 word0='d122248;
#10 word0='d122285;
#10 word0='d122322;
#10 word0='d122359;
#10 word0='d122396;
#10 word0='d122433;
#10 word0='d122470;
#10 word0='d122507;
#10 word0='d122544;
#10 word0='d122581;
#10 word0='d122618;
#10 word0='d122655;
#10 word0='d122692;
#10 word0='d122729;
#10 word0='d122766;
#10 word0='d122803;
#10 word0='d122840;
#10 word0='d122877;
#10 word0='d122914;
#10 word0='d122951;
#10 word0='d122988;
#10 word0='d123025;
#10 word0='d123062;
#10 word0='d123099;
#10 word0='d123136;
#10 word0='d123173;
#10 word0='d123210;
#10 word0='d123247;
#10 word0='d123284;
#10 word0='d123321;
#10 word0='d123358;
#10 word0='d123395;
#10 word0='d123432;
#10 word0='d123469;
#10 word0='d123506;
#10 word0='d123543;
#10 word0='d123580;
#10 word0='d123617;
#10 word0='d123654;
#10 word0='d123691;
#10 word0='d123728;
#10 word0='d123765;
#10 word0='d123802;
#10 word0='d123839;
#10 word0='d123876;
#10 word0='d123913;
#10 word0='d123950;
#10 word0='d123987;
#10 word0='d124024;
#10 word0='d124061;
#10 word0='d124098;
#10 word0='d124135;
#10 word0='d124172;
#10 word0='d124209;
#10 word0='d124246;
#10 word0='d124283;
#10 word0='d124320;
#10 word0='d124357;
#10 word0='d124394;
#10 word0='d124431;
#10 word0='d124468;
#10 word0='d124505;
#10 word0='d124542;
#10 word0='d124579;
#10 word0='d124616;
#10 word0='d124653;
#10 word0='d124690;
#10 word0='d124727;
#10 word0='d124764;
#10 word0='d124801;
#10 word0='d124838;
#10 word0='d124875;
#10 word0='d124912;
#10 word0='d124949;
#10 word0='d124986;
#10 word0='d125023;
#10 word0='d125060;
#10 word0='d125097;
#10 word0='d125134;
#10 word0='d125171;
#10 word0='d125208;
#10 word0='d125245;
#10 word0='d125282;
#10 word0='d125319;
#10 word0='d125356;
#10 word0='d125393;
#10 word0='d125430;
#10 word0='d125467;
#10 word0='d125504;
#10 word0='d125541;
#10 word0='d125578;
#10 word0='d125615;
#10 word0='d125652;
#10 word0='d125689;
#10 word0='d125726;
#10 word0='d125763;
#10 word0='d125800;
#10 word0='d125837;
#10 word0='d125874;
#10 word0='d125911;
#10 word0='d125948;
#10 word0='d125985;
#10 word0='d126022;
#10 word0='d126059;
#10 word0='d126096;
#10 word0='d126133;
#10 word0='d126170;
#10 word0='d126207;
#10 word0='d126244;
#10 word0='d126281;
#10 word0='d126318;
#10 word0='d126355;
#10 word0='d126392;
#10 word0='d126429;
#10 word0='d126466;
#10 word0='d126503;
#10 word0='d126540;
#10 word0='d126577;
#10 word0='d126614;
#10 word0='d126651;
#10 word0='d126688;
#10 word0='d126725;
#10 word0='d126762;
#10 word0='d126799;
#10 word0='d126836;
#10 word0='d126873;
#10 word0='d126910;
#10 word0='d126947;
#10 word0='d126984;
#10 word0='d127021;
#10 word0='d127058;
#10 word0='d127095;
#10 word0='d127132;
#10 word0='d127169;
#10 word0='d127206;
#10 word0='d127243;
#10 word0='d127280;
#10 word0='d127317;
#10 word0='d127354;
#10 word0='d127391;
#10 word0='d127428;
#10 word0='d127465;
#10 word0='d127502;
#10 word0='d127539;
#10 word0='d127576;
#10 word0='d127613;
#10 word0='d127650;
#10 word0='d127687;
#10 word0='d127724;
#10 word0='d127761;
#10 word0='d127798;
#10 word0='d127835;
#10 word0='d127872;
#10 word0='d127909;
#10 word0='d127946;
#10 word0='d127983;
#10 word0='d128020;
#10 word0='d128057;
#10 word0='d128094;
#10 word0='d128131;
#10 word0='d128168;
#10 word0='d128205;
#10 word0='d128242;
#10 word0='d128279;
#10 word0='d128316;
#10 word0='d128353;
#10 word0='d128390;
#10 word0='d128427;
#10 word0='d128464;
#10 word0='d128501;
#10 word0='d128538;
#10 word0='d128575;
#10 word0='d128612;
#10 word0='d128649;
#10 word0='d128686;
#10 word0='d128723;
#10 word0='d128760;
#10 word0='d128797;
#10 word0='d128834;
#10 word0='d128871;
#10 word0='d128908;
#10 word0='d128945;
#10 word0='d128982;
#10 word0='d129019;
#10 word0='d129056;
#10 word0='d129093;
#10 word0='d129130;
#10 word0='d129167;
#10 word0='d129204;
#10 word0='d129241;
#10 word0='d129278;
#10 word0='d129315;
#10 word0='d129352;
#10 word0='d129389;
#10 word0='d129426;
#10 word0='d129463;
#10 word0='d129500;
#10 word0='d129537;
#10 word0='d129574;
#10 word0='d129611;
#10 word0='d129648;
#10 word0='d129685;
#10 word0='d129722;
#10 word0='d129759;
#10 word0='d129796;
#10 word0='d129833;
#10 word0='d129870;
#10 word0='d129907;
#10 word0='d129944;
#10 word0='d129981;
#10 word0='d130018;
#10 word0='d130055;
#10 word0='d130092;
#10 word0='d130129;
#10 word0='d130166;
#10 word0='d130203;
#10 word0='d130240;
#10 word0='d130277;
#10 word0='d130314;
#10 word0='d130351;
#10 word0='d130388;
#10 word0='d130425;
#10 word0='d130462;
#10 word0='d130499;
#10 word0='d130536;
#10 word0='d130573;
#10 word0='d130610;
#10 word0='d130647;
#10 word0='d130684;
#10 word0='d130721;
#10 word0='d130758;
#10 word0='d130795;
#10 word0='d130832;
#10 word0='d130869;
#10 word0='d130906;
#10 word0='d130943;
#10 word0='d130980;
#10 word0='d131017;
#10 word0='d131054;
#10 word0='d131091;
#10 word0='d131128;
#10 word0='d131165;
#10 word0='d131202;
#10 word0='d131239;
#10 word0='d131276;
#10 word0='d131313;
#10 word0='d131350;
#10 word0='d131387;
#10 word0='d131424;
#10 word0='d131461;
#10 word0='d131498;
#10 word0='d131535;
#10 word0='d131572;
#10 word0='d131609;
#10 word0='d131646;
#10 word0='d131683;
#10 word0='d131720;
#10 word0='d131757;
#10 word0='d131794;
#10 word0='d131831;
#10 word0='d131868;
#10 word0='d131905;
#10 word0='d131942;
#10 word0='d131979;
#10 word0='d132016;
#10 word0='d132053;
#10 word0='d132090;
#10 word0='d132127;
#10 word0='d132164;
#10 word0='d132201;
#10 word0='d132238;
#10 word0='d132275;
#10 word0='d132312;
#10 word0='d132349;
#10 word0='d132386;
#10 word0='d132423;
#10 word0='d132460;
#10 word0='d132497;
#10 word0='d132534;
#10 word0='d132571;
#10 word0='d132608;
#10 word0='d132645;
#10 word0='d132682;
#10 word0='d132719;
#10 word0='d132756;
#10 word0='d132793;
#10 word0='d132830;
#10 word0='d132867;
#10 word0='d132904;
#10 word0='d132941;
#10 word0='d132978;
#10 word0='d133015;
#10 word0='d133052;
#10 word0='d133089;
#10 word0='d133126;
#10 word0='d133163;
#10 word0='d133200;
#10 word0='d133237;
#10 word0='d133274;
#10 word0='d133311;
#10 word0='d133348;
#10 word0='d133385;
#10 word0='d133422;
#10 word0='d133459;
#10 word0='d133496;
#10 word0='d133533;
#10 word0='d133570;
#10 word0='d133607;
#10 word0='d133644;
#10 word0='d133681;
#10 word0='d133718;
#10 word0='d133755;
#10 word0='d133792;
#10 word0='d133829;
#10 word0='d133866;
#10 word0='d133903;
#10 word0='d133940;
#10 word0='d133977;
#10 word0='d134014;
#10 word0='d134051;
#10 word0='d134088;
#10 word0='d134125;
#10 word0='d134162;
#10 word0='d134199;
#10 word0='d134236;
#10 word0='d134273;
#10 word0='d134310;
#10 word0='d134347;
#10 word0='d134384;
#10 word0='d134421;
#10 word0='d134458;
#10 word0='d134495;
#10 word0='d134532;
#10 word0='d134569;
#10 word0='d134606;
#10 word0='d134643;
#10 word0='d134680;
#10 word0='d134717;
#10 word0='d134754;
#10 word0='d134791;
#10 word0='d134828;
#10 word0='d134865;
#10 word0='d134902;
#10 word0='d134939;
#10 word0='d134976;
#10 word0='d135013;
#10 word0='d135050;
#10 word0='d135087;
#10 word0='d135124;
#10 word0='d135161;
#10 word0='d135198;
#10 word0='d135235;
#10 word0='d135272;
#10 word0='d135309;
#10 word0='d135346;
#10 word0='d135383;
#10 word0='d135420;
#10 word0='d135457;
#10 word0='d135494;
#10 word0='d135531;
#10 word0='d135568;
#10 word0='d135605;
#10 word0='d135642;
#10 word0='d135679;
#10 word0='d135716;
#10 word0='d135753;
#10 word0='d135790;
#10 word0='d135827;
#10 word0='d135864;
#10 word0='d135901;
#10 word0='d135938;
#10 word0='d135975;
#10 word0='d136012;
#10 word0='d136049;
#10 word0='d136086;
#10 word0='d136123;
#10 word0='d136160;
#10 word0='d136197;
#10 word0='d136234;
#10 word0='d136271;
#10 word0='d136308;
#10 word0='d136345;
#10 word0='d136382;
#10 word0='d136419;
#10 word0='d136456;
#10 word0='d136493;
#10 word0='d136530;
#10 word0='d136567;
#10 word0='d136604;
#10 word0='d136641;
#10 word0='d136678;
#10 word0='d136715;
#10 word0='d136752;
#10 word0='d136789;
#10 word0='d136826;
#10 word0='d136863;
#10 word0='d136900;
#10 word0='d136937;
#10 word0='d136974;
#10 word0='d137011;
#10 word0='d137048;
#10 word0='d137085;
#10 word0='d137122;
#10 word0='d137159;
#10 word0='d137196;
#10 word0='d137233;
#10 word0='d137270;
#10 word0='d137307;
#10 word0='d137344;
#10 word0='d137381;
#10 word0='d137418;
#10 word0='d137455;
#10 word0='d137492;
#10 word0='d137529;
#10 word0='d137566;
#10 word0='d137603;
#10 word0='d137640;
#10 word0='d137677;
#10 word0='d137714;
#10 word0='d137751;
#10 word0='d137788;
#10 word0='d137825;
#10 word0='d137862;
#10 word0='d137899;
#10 word0='d137936;
#10 word0='d137973;
#10 word0='d138010;
#10 word0='d138047;
#10 word0='d138084;
#10 word0='d138121;
#10 word0='d138158;
#10 word0='d138195;
#10 word0='d138232;
#10 word0='d138269;
#10 word0='d138306;
#10 word0='d138343;
#10 word0='d138380;
#10 word0='d138417;
#10 word0='d138454;
#10 word0='d138491;
#10 word0='d138528;
#10 word0='d138565;
#10 word0='d138602;
#10 word0='d138639;
#10 word0='d138676;
#10 word0='d138713;
#10 word0='d138750;
#10 word0='d138787;
#10 word0='d138824;
#10 word0='d138861;
#10 word0='d138898;
#10 word0='d138935;
#10 word0='d138972;
#10 word0='d139009;
#10 word0='d139046;
#10 word0='d139083;
#10 word0='d139120;
#10 word0='d139157;
#10 word0='d139194;
#10 word0='d139231;
#10 word0='d139268;
#10 word0='d139305;
#10 word0='d139342;
#10 word0='d139379;
#10 word0='d139416;
#10 word0='d139453;
#10 word0='d139490;
#10 word0='d139527;
#10 word0='d139564;
#10 word0='d139601;
#10 word0='d139638;
#10 word0='d139675;
#10 word0='d139712;
#10 word0='d139749;
#10 word0='d139786;
#10 word0='d139823;
#10 word0='d139860;
#10 word0='d139897;
#10 word0='d139934;
#10 word0='d139971;
#10 word0='d140008;
#10 word0='d140045;
#10 word0='d140082;
#10 word0='d140119;
#10 word0='d140156;
#10 word0='d140193;
#10 word0='d140230;
#10 word0='d140267;
#10 word0='d140304;
#10 word0='d140341;
#10 word0='d140378;
#10 word0='d140415;
#10 word0='d140452;
#10 word0='d140489;
#10 word0='d140526;
#10 word0='d140563;
#10 word0='d140600;
#10 word0='d140637;
#10 word0='d140674;
#10 word0='d140711;
#10 word0='d140748;
#10 word0='d140785;
#10 word0='d140822;
#10 word0='d140859;
#10 word0='d140896;
#10 word0='d140933;
#10 word0='d140970;
#10 word0='d141007;
#10 word0='d141044;
#10 word0='d141081;
#10 word0='d141118;
#10 word0='d141155;
#10 word0='d141192;
#10 word0='d141229;
#10 word0='d141266;
#10 word0='d141303;
#10 word0='d141340;
#10 word0='d141377;
#10 word0='d141414;
#10 word0='d141451;
#10 word0='d141488;
#10 word0='d141525;
#10 word0='d141562;
#10 word0='d141599;
#10 word0='d141636;
#10 word0='d141673;
#10 word0='d141710;
#10 word0='d141747;
#10 word0='d141784;
#10 word0='d141821;
#10 word0='d141858;
#10 word0='d141895;
#10 word0='d141932;
#10 word0='d141969;
#10 word0='d142006;
#10 word0='d142043;
#10 word0='d142080;
#10 word0='d142117;
#10 word0='d142154;
#10 word0='d142191;
#10 word0='d142228;
#10 word0='d142265;
#10 word0='d142302;
#10 word0='d142339;
#10 word0='d142376;
#10 word0='d142413;
#10 word0='d142450;
#10 word0='d142487;
#10 word0='d142524;
#10 word0='d142561;
#10 word0='d142598;
#10 word0='d142635;
#10 word0='d142672;
#10 word0='d142709;
#10 word0='d142746;
#10 word0='d142783;
#10 word0='d142820;
#10 word0='d142857;
#10 word0='d142894;
#10 word0='d142931;
#10 word0='d142968;
#10 word0='d143005;
#10 word0='d143042;
#10 word0='d143079;
#10 word0='d143116;
#10 word0='d143153;
#10 word0='d143190;
#10 word0='d143227;
#10 word0='d143264;
#10 word0='d143301;
#10 word0='d143338;
#10 word0='d143375;
#10 word0='d143412;
#10 word0='d143449;
#10 word0='d143486;
#10 word0='d143523;
#10 word0='d143560;
#10 word0='d143597;
#10 word0='d143634;
#10 word0='d143671;
#10 word0='d143708;
#10 word0='d143745;
#10 word0='d143782;
#10 word0='d143819;
#10 word0='d143856;
#10 word0='d143893;
#10 word0='d143930;
#10 word0='d143967;
#10 word0='d144004;
#10 word0='d144041;
#10 word0='d144078;
#10 word0='d144115;
#10 word0='d144152;
#10 word0='d144189;
#10 word0='d144226;
#10 word0='d144263;
#10 word0='d144300;
#10 word0='d144337;
#10 word0='d144374;
#10 word0='d144411;
#10 word0='d144448;
#10 word0='d144485;
#10 word0='d144522;
#10 word0='d144559;
#10 word0='d144596;
#10 word0='d144633;
#10 word0='d144670;
#10 word0='d144707;
#10 word0='d144744;
#10 word0='d144781;
#10 word0='d144818;
#10 word0='d144855;
#10 word0='d144892;
#10 word0='d144929;
#10 word0='d144966;
#10 word0='d145003;
#10 word0='d145040;
#10 word0='d145077;
#10 word0='d145114;
#10 word0='d145151;
#10 word0='d145188;
#10 word0='d145225;
#10 word0='d145262;
#10 word0='d145299;
#10 word0='d145336;
#10 word0='d145373;
#10 word0='d145410;
#10 word0='d145447;
#10 word0='d145484;
#10 word0='d145521;
#10 word0='d145558;
#10 word0='d145595;
#10 word0='d145632;
#10 word0='d145669;
#10 word0='d145706;
#10 word0='d145743;
#10 word0='d145780;
#10 word0='d145817;
#10 word0='d145854;
#10 word0='d145891;
#10 word0='d145928;
#10 word0='d145965;
#10 word0='d146002;
#10 word0='d146039;
#10 word0='d146076;
#10 word0='d146113;
#10 word0='d146150;
#10 word0='d146187;
#10 word0='d146224;
#10 word0='d146261;
#10 word0='d146298;
#10 word0='d146335;
#10 word0='d146372;
#10 word0='d146409;
#10 word0='d146446;
#10 word0='d146483;
#10 word0='d146520;
#10 word0='d146557;
#10 word0='d146594;
#10 word0='d146631;
#10 word0='d146668;
#10 word0='d146705;
#10 word0='d146742;
#10 word0='d146779;
#10 word0='d146816;
#10 word0='d146853;
#10 word0='d146890;
#10 word0='d146927;
#10 word0='d146964;
#10 word0='d147001;
#10 word0='d147038;
#10 word0='d147075;
#10 word0='d147112;
#10 word0='d147149;
#10 word0='d147186;
#10 word0='d147223;
#10 word0='d147260;
#10 word0='d147297;
#10 word0='d147334;
#10 word0='d147371;
#10 word0='d147408;
#10 word0='d147445;
#10 word0='d147482;
#10 word0='d147519;
#10 word0='d147556;
#10 word0='d147593;
#10 word0='d147630;
#10 word0='d147667;
#10 word0='d147704;
#10 word0='d147741;
#10 word0='d147778;
#10 word0='d147815;
#10 word0='d147852;
#10 word0='d147889;
#10 word0='d147926;
#10 word0='d147963;
#10 word0='d148000;
#10 word0='d148037;
#10 word0='d148074;
#10 word0='d148111;
#10 word0='d148148;
#10 word0='d148185;
#10 word0='d148222;
#10 word0='d148259;
#10 word0='d148296;
#10 word0='d148333;
#10 word0='d148370;
#10 word0='d148407;
#10 word0='d148444;
#10 word0='d148481;
#10 word0='d148518;
#10 word0='d148555;
#10 word0='d148592;
#10 word0='d148629;
#10 word0='d148666;
#10 word0='d148703;
#10 word0='d148740;
#10 word0='d148777;
#10 word0='d148814;
#10 word0='d148851;
#10 word0='d148888;
#10 word0='d148925;
#10 word0='d148962;
#10 word0='d148999;
#10 word0='d149036;
#10 word0='d149073;
#10 word0='d149110;
#10 word0='d149147;
#10 word0='d149184;
#10 word0='d149221;
#10 word0='d149258;
#10 word0='d149295;
#10 word0='d149332;
#10 word0='d149369;
#10 word0='d149406;
#10 word0='d149443;
#10 word0='d149480;
#10 word0='d149517;
#10 word0='d149554;
#10 word0='d149591;
#10 word0='d149628;
#10 word0='d149665;
#10 word0='d149702;
#10 word0='d149739;
#10 word0='d149776;
#10 word0='d149813;
#10 word0='d149850;
#10 word0='d149887;
#10 word0='d149924;
#10 word0='d149961;
#10 word0='d149998;
#10 word0='d150035;
#10 word0='d150072;
#10 word0='d150109;
#10 word0='d150146;
#10 word0='d150183;
#10 word0='d150220;
#10 word0='d150257;
#10 word0='d150294;
#10 word0='d150331;
#10 word0='d150368;
#10 word0='d150405;
#10 word0='d150442;
#10 word0='d150479;
#10 word0='d150516;
#10 word0='d150553;
#10 word0='d150590;
#10 word0='d150627;
#10 word0='d150664;
#10 word0='d150701;
#10 word0='d150738;
#10 word0='d150775;
#10 word0='d150812;
#10 word0='d150849;
#10 word0='d150886;
#10 word0='d150923;
#10 word0='d150960;
#10 word0='d150997;
#10 word0='d151034;
#10 word0='d151071;
#10 word0='d151108;
#10 word0='d151145;
#10 word0='d151182;
#10 word0='d151219;
#10 word0='d151256;
#10 word0='d151293;
#10 word0='d151330;
#10 word0='d151367;
#10 word0='d151404;
#10 word0='d151441;
#10 word0='d151478;
#10 word0='d151515;
#10 word0='d151552;
#10 word0='d151589;
#10 word0='d151626;
#10 word0='d151663;
#10 word0='d151700;
#10 word0='d151737;
#10 word0='d151774;
#10 word0='d151811;
#10 word0='d151848;
#10 word0='d151885;
#10 word0='d151922;
#10 word0='d151959;
#10 word0='d151996;
#10 word0='d152033;
#10 word0='d152070;
#10 word0='d152107;
#10 word0='d152144;
#10 word0='d152181;
#10 word0='d152218;
#10 word0='d152255;
#10 word0='d152292;
#10 word0='d152329;
#10 word0='d152366;
#10 word0='d152403;
#10 word0='d152440;
#10 word0='d152477;
#10 word0='d152514;
#10 word0='d152551;
#10 word0='d152588;
#10 word0='d152625;
#10 word0='d152662;
#10 word0='d152699;
#10 word0='d152736;
#10 word0='d152773;
#10 word0='d152810;
#10 word0='d152847;
#10 word0='d152884;
#10 word0='d152921;
#10 word0='d152958;
#10 word0='d152995;
#10 word0='d153032;
#10 word0='d153069;
#10 word0='d153106;
#10 word0='d153143;
#10 word0='d153180;
#10 word0='d153217;
#10 word0='d153254;
#10 word0='d153291;
#10 word0='d153328;
#10 word0='d153365;
#10 word0='d153402;
#10 word0='d153439;
#10 word0='d153476;
#10 word0='d153513;
#10 word0='d153550;
#10 word0='d153587;
#10 word0='d153624;
#10 word0='d153661;
#10 word0='d153698;
#10 word0='d153735;
#10 word0='d153772;
#10 word0='d153809;
#10 word0='d153846;
#10 word0='d153883;
#10 word0='d153920;
#10 word0='d153957;
#10 word0='d153994;
#10 word0='d154031;
#10 word0='d154068;
#10 word0='d154105;
#10 word0='d154142;
#10 word0='d154179;
#10 word0='d154216;
#10 word0='d154253;
#10 word0='d154290;
#10 word0='d154327;
#10 word0='d154364;
#10 word0='d154401;
#10 word0='d154438;
#10 word0='d154475;
#10 word0='d154512;
#10 word0='d154549;
#10 word0='d154586;
#10 word0='d154623;
#10 word0='d154660;
#10 word0='d154697;
#10 word0='d154734;
#10 word0='d154771;
#10 word0='d154808;
#10 word0='d154845;
#10 word0='d154882;
#10 word0='d154919;
#10 word0='d154956;
#10 word0='d154993;
#10 word0='d155030;
#10 word0='d155067;
#10 word0='d155104;
#10 word0='d155141;
#10 word0='d155178;
#10 word0='d155215;
#10 word0='d155252;
#10 word0='d155289;
#10 word0='d155326;
#10 word0='d155363;
#10 word0='d155400;
#10 word0='d155437;
#10 word0='d155474;
#10 word0='d155511;
#10 word0='d155548;
#10 word0='d155585;
#10 word0='d155622;
#10 word0='d155659;
#10 word0='d155696;
#10 word0='d155733;
#10 word0='d155770;
#10 word0='d155807;
#10 word0='d155844;
#10 word0='d155881;
#10 word0='d155918;
#10 word0='d155955;
#10 word0='d155992;
#10 word0='d156029;
#10 word0='d156066;
#10 word0='d156103;
#10 word0='d156140;
#10 word0='d156177;
#10 word0='d156214;
#10 word0='d156251;
#10 word0='d156288;
#10 word0='d156325;
#10 word0='d156362;
#10 word0='d156399;
#10 word0='d156436;
#10 word0='d156473;
#10 word0='d156510;
#10 word0='d156547;
#10 word0='d156584;
#10 word0='d156621;
#10 word0='d156658;
#10 word0='d156695;
#10 word0='d156732;
#10 word0='d156769;
#10 word0='d156806;
#10 word0='d156843;
#10 word0='d156880;
#10 word0='d156917;
#10 word0='d156954;
#10 word0='d156991;
#10 word0='d157028;
#10 word0='d157065;
#10 word0='d157102;
#10 word0='d157139;
#10 word0='d157176;
#10 word0='d157213;
#10 word0='d157250;
#10 word0='d157287;
#10 word0='d157324;
#10 word0='d157361;
#10 word0='d157398;
#10 word0='d157435;
#10 word0='d157472;
#10 word0='d157509;
#10 word0='d157546;
#10 word0='d157583;
#10 word0='d157620;
#10 word0='d157657;
#10 word0='d157694;
#10 word0='d157731;
#10 word0='d157768;
#10 word0='d157805;
#10 word0='d157842;
#10 word0='d157879;
#10 word0='d157916;
#10 word0='d157953;
#10 word0='d157990;
#10 word0='d158027;
#10 word0='d158064;
#10 word0='d158101;
#10 word0='d158138;
#10 word0='d158175;
#10 word0='d158212;
#10 word0='d158249;
#10 word0='d158286;
#10 word0='d158323;
#10 word0='d158360;
#10 word0='d158397;
#10 word0='d158434;
#10 word0='d158471;
#10 word0='d158508;
#10 word0='d158545;
#10 word0='d158582;
#10 word0='d158619;
#10 word0='d158656;
#10 word0='d158693;
#10 word0='d158730;
#10 word0='d158767;
#10 word0='d158804;
#10 word0='d158841;
#10 word0='d158878;
#10 word0='d158915;
#10 word0='d158952;
#10 word0='d158989;
#10 word0='d159026;
#10 word0='d159063;
#10 word0='d159100;
#10 word0='d159137;
#10 word0='d159174;
#10 word0='d159211;
#10 word0='d159248;
#10 word0='d159285;
#10 word0='d159322;
#10 word0='d159359;
#10 word0='d159396;
#10 word0='d159433;
#10 word0='d159470;
#10 word0='d159507;
#10 word0='d159544;
#10 word0='d159581;
#10 word0='d159618;
#10 word0='d159655;
#10 word0='d159692;
#10 word0='d159729;
#10 word0='d159766;
#10 word0='d159803;
#10 word0='d159840;
#10 word0='d159877;
#10 word0='d159914;
#10 word0='d159951;
#10 word0='d159988;
#10 word0='d160025;
#10 word0='d160062;
#10 word0='d160099;
#10 word0='d160136;
#10 word0='d160173;
#10 word0='d160210;
#10 word0='d160247;
#10 word0='d160284;
#10 word0='d160321;
#10 word0='d160358;
#10 word0='d160395;
#10 word0='d160432;
#10 word0='d160469;
#10 word0='d160506;
#10 word0='d160543;
#10 word0='d160580;
#10 word0='d160617;
#10 word0='d160654;
#10 word0='d160691;
#10 word0='d160728;
#10 word0='d160765;
#10 word0='d160802;
#10 word0='d160839;
#10 word0='d160876;
#10 word0='d160913;
#10 word0='d160950;
#10 word0='d160987;
#10 word0='d161024;
#10 word0='d161061;
#10 word0='d161098;
#10 word0='d161135;
#10 word0='d161172;
#10 word0='d161209;
#10 word0='d161246;
#10 word0='d161283;
#10 word0='d161320;
#10 word0='d161357;
#10 word0='d161394;
#10 word0='d161431;
#10 word0='d161468;
#10 word0='d161505;
#10 word0='d161542;
#10 word0='d161579;
#10 word0='d161616;
#10 word0='d161653;
#10 word0='d161690;
#10 word0='d161727;
#10 word0='d161764;
#10 word0='d161801;
#10 word0='d161838;
#10 word0='d161875;
#10 word0='d161912;
#10 word0='d161949;
#10 word0='d161986;
#10 word0='d162023;
#10 word0='d162060;
#10 word0='d162097;
#10 word0='d162134;
#10 word0='d162171;
#10 word0='d162208;
#10 word0='d162245;
#10 word0='d162282;
#10 word0='d162319;
#10 word0='d162356;
#10 word0='d162393;
#10 word0='d162430;
#10 word0='d162467;
#10 word0='d162504;
#10 word0='d162541;
#10 word0='d162578;
#10 word0='d162615;
#10 word0='d162652;
#10 word0='d162689;
#10 word0='d162726;
#10 word0='d162763;
#10 word0='d162800;
#10 word0='d162837;
#10 word0='d162874;
#10 word0='d162911;
#10 word0='d162948;
#10 word0='d162985;
#10 word0='d163022;
#10 word0='d163059;
#10 word0='d163096;
#10 word0='d163133;
#10 word0='d163170;
#10 word0='d163207;
#10 word0='d163244;
#10 word0='d163281;
#10 word0='d163318;
#10 word0='d163355;
#10 word0='d163392;
#10 word0='d163429;
#10 word0='d163466;
#10 word0='d163503;
#10 word0='d163540;
#10 word0='d163577;
#10 word0='d163614;
#10 word0='d163651;
#10 word0='d163688;
#10 word0='d163725;
#10 word0='d163762;
#10 word0='d163799;
#10 word0='d163836;
#10 word0='d163873;
#10 word0='d163910;
#10 word0='d163947;
#10 word0='d163984;
#10 word0='d164021;
#10 word0='d164058;
#10 word0='d164095;
#10 word0='d164132;
#10 word0='d164169;
#10 word0='d164206;
#10 word0='d164243;
#10 word0='d164280;
#10 word0='d164317;
#10 word0='d164354;
#10 word0='d164391;
#10 word0='d164428;
#10 word0='d164465;
#10 word0='d164502;
#10 word0='d164539;
#10 word0='d164576;
#10 word0='d164613;
#10 word0='d164650;
#10 word0='d164687;
#10 word0='d164724;
#10 word0='d164761;
#10 word0='d164798;
#10 word0='d164835;
#10 word0='d164872;
#10 word0='d164909;
#10 word0='d164946;
#10 word0='d164983;
#10 word0='d165020;
#10 word0='d165057;
#10 word0='d165094;
#10 word0='d165131;
#10 word0='d165168;
#10 word0='d165205;
#10 word0='d165242;
#10 word0='d165279;
#10 word0='d165316;
#10 word0='d165353;
#10 word0='d165390;
#10 word0='d165427;
#10 word0='d165464;
#10 word0='d165501;
#10 word0='d165538;
#10 word0='d165575;
#10 word0='d165612;
#10 word0='d165649;
#10 word0='d165686;
#10 word0='d165723;
#10 word0='d165760;
#10 word0='d165797;
#10 word0='d165834;
#10 word0='d165871;
#10 word0='d165908;
#10 word0='d165945;
#10 word0='d165982;
#10 word0='d166019;
#10 word0='d166056;
#10 word0='d166093;
#10 word0='d166130;
#10 word0='d166167;
#10 word0='d166204;
#10 word0='d166241;
#10 word0='d166278;
#10 word0='d166315;
#10 word0='d166352;
#10 word0='d166389;
#10 word0='d166426;
#10 word0='d166463;
#10 word0='d166500;
#10 word0='d166537;
#10 word0='d166574;
#10 word0='d166611;
#10 word0='d166648;
#10 word0='d166685;
#10 word0='d166722;
#10 word0='d166759;
#10 word0='d166796;
#10 word0='d166833;
#10 word0='d166870;
#10 word0='d166907;
#10 word0='d166944;
#10 word0='d166981;
#10 word0='d167018;
#10 word0='d167055;
#10 word0='d167092;
#10 word0='d167129;
#10 word0='d167166;
#10 word0='d167203;
#10 word0='d167240;
#10 word0='d167277;
#10 word0='d167314;
#10 word0='d167351;
#10 word0='d167388;
#10 word0='d167425;
#10 word0='d167462;
#10 word0='d167499;
#10 word0='d167536;
#10 word0='d167573;
#10 word0='d167610;
#10 word0='d167647;
#10 word0='d167684;
#10 word0='d167721;
#10 word0='d167758;
#10 word0='d167795;
#10 word0='d167832;
#10 word0='d167869;
#10 word0='d167906;
#10 word0='d167943;
#10 word0='d167980;
#10 word0='d168017;
#10 word0='d168054;
#10 word0='d168091;
#10 word0='d168128;
#10 word0='d168165;
#10 word0='d168202;
#10 word0='d168239;
#10 word0='d168276;
#10 word0='d168313;
#10 word0='d168350;
#10 word0='d168387;
#10 word0='d168424;
#10 word0='d168461;
#10 word0='d168498;
#10 word0='d168535;
#10 word0='d168572;
#10 word0='d168609;
#10 word0='d168646;
#10 word0='d168683;
#10 word0='d168720;
#10 word0='d168757;
#10 word0='d168794;
#10 word0='d168831;
#10 word0='d168868;
#10 word0='d168905;
#10 word0='d168942;
#10 word0='d168979;
#10 word0='d169016;
#10 word0='d169053;
#10 word0='d169090;
#10 word0='d169127;
#10 word0='d169164;
#10 word0='d169201;
#10 word0='d169238;
#10 word0='d169275;
#10 word0='d169312;
#10 word0='d169349;
#10 word0='d169386;
#10 word0='d169423;
#10 word0='d169460;
#10 word0='d169497;
#10 word0='d169534;
#10 word0='d169571;
#10 word0='d169608;
#10 word0='d169645;
#10 word0='d169682;
#10 word0='d169719;
#10 word0='d169756;
#10 word0='d169793;
#10 word0='d169830;
#10 word0='d169867;
#10 word0='d169904;
#10 word0='d169941;
#10 word0='d169978;
#10 word0='d170015;
#10 word0='d170052;
#10 word0='d170089;
#10 word0='d170126;
#10 word0='d170163;
#10 word0='d170200;
#10 word0='d170237;
#10 word0='d170274;
#10 word0='d170311;
#10 word0='d170348;
#10 word0='d170385;
#10 word0='d170422;
#10 word0='d170459;
#10 word0='d170496;
#10 word0='d170533;
#10 word0='d170570;
#10 word0='d170607;
#10 word0='d170644;
#10 word0='d170681;
#10 word0='d170718;
#10 word0='d170755;
#10 word0='d170792;
#10 word0='d170829;
#10 word0='d170866;
#10 word0='d170903;
#10 word0='d170940;
#10 word0='d170977;
#10 word0='d171014;
#10 word0='d171051;
#10 word0='d171088;
#10 word0='d171125;
#10 word0='d171162;
#10 word0='d171199;
#10 word0='d171236;
#10 word0='d171273;
#10 word0='d171310;
#10 word0='d171347;
#10 word0='d171384;
#10 word0='d171421;
#10 word0='d171458;
#10 word0='d171495;
#10 word0='d171532;
#10 word0='d171569;
#10 word0='d171606;
#10 word0='d171643;
#10 word0='d171680;
#10 word0='d171717;
#10 word0='d171754;
#10 word0='d171791;
#10 word0='d171828;
#10 word0='d171865;
#10 word0='d171902;
#10 word0='d171939;
#10 word0='d171976;
#10 word0='d172013;
#10 word0='d172050;
#10 word0='d172087;
#10 word0='d172124;
#10 word0='d172161;
#10 word0='d172198;
#10 word0='d172235;
#10 word0='d172272;
#10 word0='d172309;
#10 word0='d172346;
#10 word0='d172383;
#10 word0='d172420;
#10 word0='d172457;
#10 word0='d172494;
#10 word0='d172531;
#10 word0='d172568;
#10 word0='d172605;
#10 word0='d172642;
#10 word0='d172679;
#10 word0='d172716;
#10 word0='d172753;
#10 word0='d172790;
#10 word0='d172827;
#10 word0='d172864;
#10 word0='d172901;
#10 word0='d172938;
#10 word0='d172975;
#10 word0='d173012;
#10 word0='d173049;
#10 word0='d173086;
#10 word0='d173123;
#10 word0='d173160;
#10 word0='d173197;
#10 word0='d173234;
#10 word0='d173271;
#10 word0='d173308;
#10 word0='d173345;
#10 word0='d173382;
#10 word0='d173419;
#10 word0='d173456;
#10 word0='d173493;
#10 word0='d173530;
#10 word0='d173567;
#10 word0='d173604;
#10 word0='d173641;
#10 word0='d173678;
#10 word0='d173715;
#10 word0='d173752;
#10 word0='d173789;
#10 word0='d173826;
#10 word0='d173863;
#10 word0='d173900;
#10 word0='d173937;
#10 word0='d173974;
#10 word0='d174011;
#10 word0='d174048;
#10 word0='d174085;
#10 word0='d174122;
#10 word0='d174159;
#10 word0='d174196;
#10 word0='d174233;
#10 word0='d174270;
#10 word0='d174307;
#10 word0='d174344;
#10 word0='d174381;
#10 word0='d174418;
#10 word0='d174455;
#10 word0='d174492;
#10 word0='d174529;
#10 word0='d174566;
#10 word0='d174603;
#10 word0='d174640;
#10 word0='d174677;
#10 word0='d174714;
#10 word0='d174751;
#10 word0='d174788;
#10 word0='d174825;
#10 word0='d174862;
#10 word0='d174899;
#10 word0='d174936;
#10 word0='d174973;
#10 word0='d175010;
#10 word0='d175047;
#10 word0='d175084;
#10 word0='d175121;
#10 word0='d175158;
#10 word0='d175195;
#10 word0='d175232;
#10 word0='d175269;
#10 word0='d175306;
#10 word0='d175343;
#10 word0='d175380;
#10 word0='d175417;
#10 word0='d175454;
#10 word0='d175491;
#10 word0='d175528;
#10 word0='d175565;
#10 word0='d175602;
#10 word0='d175639;
#10 word0='d175676;
#10 word0='d175713;
#10 word0='d175750;
#10 word0='d175787;
#10 word0='d175824;
#10 word0='d175861;
#10 word0='d175898;
#10 word0='d175935;
#10 word0='d175972;
#10 word0='d176009;
#10 word0='d176046;
#10 word0='d176083;
#10 word0='d176120;
#10 word0='d176157;
#10 word0='d176194;
#10 word0='d176231;
#10 word0='d176268;
#10 word0='d176305;
#10 word0='d176342;
#10 word0='d176379;
#10 word0='d176416;
#10 word0='d176453;
#10 word0='d176490;
#10 word0='d176527;
#10 word0='d176564;
#10 word0='d176601;
#10 word0='d176638;
#10 word0='d176675;
#10 word0='d176712;
#10 word0='d176749;
#10 word0='d176786;
#10 word0='d176823;
#10 word0='d176860;
#10 word0='d176897;
#10 word0='d176934;
#10 word0='d176971;
#10 word0='d177008;
#10 word0='d177045;
#10 word0='d177082;
#10 word0='d177119;
#10 word0='d177156;
#10 word0='d177193;
#10 word0='d177230;
#10 word0='d177267;
#10 word0='d177304;
#10 word0='d177341;
#10 word0='d177378;
#10 word0='d177415;
#10 word0='d177452;
#10 word0='d177489;
#10 word0='d177526;
#10 word0='d177563;
#10 word0='d177600;
#10 word0='d177637;
#10 word0='d177674;
#10 word0='d177711;
#10 word0='d177748;
#10 word0='d177785;
#10 word0='d177822;
#10 word0='d177859;
#10 word0='d177896;
#10 word0='d177933;
#10 word0='d177970;
#10 word0='d178007;
#10 word0='d178044;
#10 word0='d178081;
#10 word0='d178118;
#10 word0='d178155;
#10 word0='d178192;
#10 word0='d178229;
#10 word0='d178266;
#10 word0='d178303;
#10 word0='d178340;
#10 word0='d178377;
#10 word0='d178414;
#10 word0='d178451;
#10 word0='d178488;
#10 word0='d178525;
#10 word0='d178562;
#10 word0='d178599;
#10 word0='d178636;
#10 word0='d178673;
#10 word0='d178710;
#10 word0='d178747;
#10 word0='d178784;
#10 word0='d178821;
#10 word0='d178858;
#10 word0='d178895;
#10 word0='d178932;
#10 word0='d178969;
#10 word0='d179006;
#10 word0='d179043;
#10 word0='d179080;
#10 word0='d179117;
#10 word0='d179154;
#10 word0='d179191;
#10 word0='d179228;
#10 word0='d179265;
#10 word0='d179302;
#10 word0='d179339;
#10 word0='d179376;
#10 word0='d179413;
#10 word0='d179450;
#10 word0='d179487;
#10 word0='d179524;
#10 word0='d179561;
#10 word0='d179598;
#10 word0='d179635;
#10 word0='d179672;
#10 word0='d179709;
#10 word0='d179746;
#10 word0='d179783;
#10 word0='d179820;
#10 word0='d179857;
#10 word0='d179894;
#10 word0='d179931;
#10 word0='d179968;
#10 word0='d180005;
#10 word0='d180042;
#10 word0='d180079;
#10 word0='d180116;
#10 word0='d180153;
#10 word0='d180190;
#10 word0='d180227;
#10 word0='d180264;
#10 word0='d180301;
#10 word0='d180338;
#10 word0='d180375;
#10 word0='d180412;
#10 word0='d180449;
#10 word0='d180486;
#10 word0='d180523;
#10 word0='d180560;
#10 word0='d180597;
#10 word0='d180634;
#10 word0='d180671;
#10 word0='d180708;
#10 word0='d180745;
#10 word0='d180782;
#10 word0='d180819;
#10 word0='d180856;
#10 word0='d180893;
#10 word0='d180930;
#10 word0='d180967;
#10 word0='d181004;
#10 word0='d181041;
#10 word0='d181078;
#10 word0='d181115;
#10 word0='d181152;
#10 word0='d181189;
#10 word0='d181226;
#10 word0='d181263;
#10 word0='d181300;
#10 word0='d181337;
#10 word0='d181374;
#10 word0='d181411;
#10 word0='d181448;
#10 word0='d181485;
#10 word0='d181522;
#10 word0='d181559;
#10 word0='d181596;
#10 word0='d181633;
#10 word0='d181670;
#10 word0='d181707;
#10 word0='d181744;
#10 word0='d181781;
#10 word0='d181818;
#10 word0='d181855;
#10 word0='d181892;
#10 word0='d181929;
#10 word0='d181966;
#10 word0='d182003;
#10 word0='d182040;
#10 word0='d182077;
#10 word0='d182114;
#10 word0='d182151;
#10 word0='d182188;
#10 word0='d182225;
#10 word0='d182262;
#10 word0='d182299;
#10 word0='d182336;
#10 word0='d182373;
#10 word0='d182410;
#10 word0='d182447;
#10 word0='d182484;
#10 word0='d182521;
#10 word0='d182558;
#10 word0='d182595;
#10 word0='d182632;
#10 word0='d182669;
#10 word0='d182706;
#10 word0='d182743;
#10 word0='d182780;
#10 word0='d182817;
#10 word0='d182854;
#10 word0='d182891;
#10 word0='d182928;
#10 word0='d182965;
#10 word0='d183002;
#10 word0='d183039;
#10 word0='d183076;
#10 word0='d183113;
#10 word0='d183150;
#10 word0='d183187;
#10 word0='d183224;
#10 word0='d183261;
#10 word0='d183298;
#10 word0='d183335;
#10 word0='d183372;
#10 word0='d183409;
#10 word0='d183446;
#10 word0='d183483;
#10 word0='d183520;
#10 word0='d183557;
#10 word0='d183594;
#10 word0='d183631;
#10 word0='d183668;
#10 word0='d183705;
#10 word0='d183742;
#10 word0='d183779;
#10 word0='d183816;
#10 word0='d183853;
#10 word0='d183890;
#10 word0='d183927;
#10 word0='d183964;
#10 word0='d184001;
#10 word0='d184038;
#10 word0='d184075;
#10 word0='d184112;
#10 word0='d184149;
#10 word0='d184186;
#10 word0='d184223;
#10 word0='d184260;
#10 word0='d184297;
#10 word0='d184334;
#10 word0='d184371;
#10 word0='d184408;
#10 word0='d184445;
#10 word0='d184482;
#10 word0='d184519;
#10 word0='d184556;
#10 word0='d184593;
#10 word0='d184630;
#10 word0='d184667;
#10 word0='d184704;
#10 word0='d184741;
#10 word0='d184778;
#10 word0='d184815;
#10 word0='d184852;
#10 word0='d184889;
#10 word0='d184926;
#10 word0='d184963;
#10 word0='d185000;
#10 word0='d185037;
#10 word0='d185074;
#10 word0='d185111;
#10 word0='d185148;
#10 word0='d185185;
#10 word0='d185222;
#10 word0='d185259;
#10 word0='d185296;
#10 word0='d185333;
#10 word0='d185370;
#10 word0='d185407;
#10 word0='d185444;
#10 word0='d185481;
#10 word0='d185518;
#10 word0='d185555;
#10 word0='d185592;
#10 word0='d185629;
#10 word0='d185666;
#10 word0='d185703;
#10 word0='d185740;
#10 word0='d185777;
#10 word0='d185814;
#10 word0='d185851;
#10 word0='d185888;
#10 word0='d185925;
#10 word0='d185962;
#10 word0='d185999;
#10 word0='d186036;
#10 word0='d186073;
#10 word0='d186110;
#10 word0='d186147;
#10 word0='d186184;
#10 word0='d186221;
#10 word0='d186258;
#10 word0='d186295;
#10 word0='d186332;
#10 word0='d186369;
#10 word0='d186406;
#10 word0='d186443;
#10 word0='d186480;
#10 word0='d186517;
#10 word0='d186554;
#10 word0='d186591;
#10 word0='d186628;
#10 word0='d186665;
#10 word0='d186702;
#10 word0='d186739;
#10 word0='d186776;
#10 word0='d186813;
#10 word0='d186850;
#10 word0='d186887;
#10 word0='d186924;
#10 word0='d186961;
#10 word0='d186998;
#10 word0='d187035;
#10 word0='d187072;
#10 word0='d187109;
#10 word0='d187146;
#10 word0='d187183;
#10 word0='d187220;
#10 word0='d187257;
#10 word0='d187294;
#10 word0='d187331;
#10 word0='d187368;
#10 word0='d187405;
#10 word0='d187442;
#10 word0='d187479;
#10 word0='d187516;
#10 word0='d187553;
#10 word0='d187590;
#10 word0='d187627;
#10 word0='d187664;
#10 word0='d187701;
#10 word0='d187738;
#10 word0='d187775;
#10 word0='d187812;
#10 word0='d187849;
#10 word0='d187886;
#10 word0='d187923;
#10 word0='d187960;
#10 word0='d187997;
#10 word0='d188034;
#10 word0='d188071;
#10 word0='d188108;
#10 word0='d188145;
#10 word0='d188182;
#10 word0='d188219;
#10 word0='d188256;
#10 word0='d188293;
#10 word0='d188330;
#10 word0='d188367;
#10 word0='d188404;
#10 word0='d188441;
#10 word0='d188478;
#10 word0='d188515;
#10 word0='d188552;
#10 word0='d188589;
#10 word0='d188626;
#10 word0='d188663;
#10 word0='d188700;
#10 word0='d188737;
#10 word0='d188774;
#10 word0='d188811;
#10 word0='d188848;
#10 word0='d188885;
#10 word0='d188922;
#10 word0='d188959;
#10 word0='d188996;
#10 word0='d189033;
#10 word0='d189070;
#10 word0='d189107;
#10 word0='d189144;
#10 word0='d189181;
#10 word0='d189218;
#10 word0='d189255;
#10 word0='d189292;
#10 word0='d189329;
#10 word0='d189366;
#10 word0='d189403;
#10 word0='d189440;
#10 word0='d189477;
#10 word0='d189514;
#10 word0='d189551;
#10 word0='d189588;
#10 word0='d189625;
#10 word0='d189662;
#10 word0='d189699;
#10 word0='d189736;
#10 word0='d189773;
#10 word0='d189810;
#10 word0='d189847;
#10 word0='d189884;
#10 word0='d189921;
#10 word0='d189958;
#10 word0='d189995;
#10 word0='d190032;
#10 word0='d190069;
#10 word0='d190106;
#10 word0='d190143;
#10 word0='d190180;
#10 word0='d190217;
#10 word0='d190254;
#10 word0='d190291;
#10 word0='d190328;
#10 word0='d190365;
#10 word0='d190402;
#10 word0='d190439;
#10 word0='d190476;
#10 word0='d190513;
#10 word0='d190550;
#10 word0='d190587;
#10 word0='d190624;
#10 word0='d190661;
#10 word0='d190698;
#10 word0='d190735;
#10 word0='d190772;
#10 word0='d190809;
#10 word0='d190846;
#10 word0='d190883;
#10 word0='d190920;
#10 word0='d190957;
#10 word0='d190994;
#10 word0='d191031;
#10 word0='d191068;
#10 word0='d191105;
#10 word0='d191142;
#10 word0='d191179;
#10 word0='d191216;
#10 word0='d191253;
#10 word0='d191290;
#10 word0='d191327;
#10 word0='d191364;
#10 word0='d191401;
#10 word0='d191438;
#10 word0='d191475;
#10 word0='d191512;
#10 word0='d191549;
#10 word0='d191586;
#10 word0='d191623;
#10 word0='d191660;
#10 word0='d191697;
#10 word0='d191734;
#10 word0='d191771;
#10 word0='d191808;
#10 word0='d191845;
#10 word0='d191882;
#10 word0='d191919;
#10 word0='d191956;
#10 word0='d191993;
#10 word0='d192030;
#10 word0='d192067;
#10 word0='d192104;
#10 word0='d192141;
#10 word0='d192178;
#10 word0='d192215;
#10 word0='d192252;
#10 word0='d192289;
#10 word0='d192326;
#10 word0='d192363;
#10 word0='d192400;
#10 word0='d192437;
#10 word0='d192474;
#10 word0='d192511;
#10 word0='d192548;
#10 word0='d192585;
#10 word0='d192622;
#10 word0='d192659;
#10 word0='d192696;
#10 word0='d192733;
#10 word0='d192770;
#10 word0='d192807;
#10 word0='d192844;
#10 word0='d192881;
#10 word0='d192918;
#10 word0='d192955;
#10 word0='d192992;
#10 word0='d193029;
#10 word0='d193066;
#10 word0='d193103;
#10 word0='d193140;
#10 word0='d193177;
#10 word0='d193214;
#10 word0='d193251;
#10 word0='d193288;
#10 word0='d193325;
#10 word0='d193362;
#10 word0='d193399;
#10 word0='d193436;
#10 word0='d193473;
#10 word0='d193510;
#10 word0='d193547;
#10 word0='d193584;
#10 word0='d193621;
#10 word0='d193658;
#10 word0='d193695;
#10 word0='d193732;
#10 word0='d193769;
#10 word0='d193806;
#10 word0='d193843;
#10 word0='d193880;
#10 word0='d193917;
#10 word0='d193954;
#10 word0='d193991;
#10 word0='d194028;
#10 word0='d194065;
#10 word0='d194102;
#10 word0='d194139;
#10 word0='d194176;
#10 word0='d194213;
#10 word0='d194250;
#10 word0='d194287;
#10 word0='d194324;
#10 word0='d194361;
#10 word0='d194398;
#10 word0='d194435;
#10 word0='d194472;
#10 word0='d194509;
#10 word0='d194546;
#10 word0='d194583;
#10 word0='d194620;
#10 word0='d194657;
#10 word0='d194694;
#10 word0='d194731;
#10 word0='d194768;
#10 word0='d194805;
#10 word0='d194842;
#10 word0='d194879;
#10 word0='d194916;
#10 word0='d194953;
#10 word0='d194990;
#10 word0='d195027;
#10 word0='d195064;
#10 word0='d195101;
#10 word0='d195138;
#10 word0='d195175;
#10 word0='d195212;
#10 word0='d195249;
#10 word0='d195286;
#10 word0='d195323;
#10 word0='d195360;
#10 word0='d195397;
#10 word0='d195434;
#10 word0='d195471;
#10 word0='d195508;
#10 word0='d195545;
#10 word0='d195582;
#10 word0='d195619;
#10 word0='d195656;
#10 word0='d195693;
#10 word0='d195730;
#10 word0='d195767;
#10 word0='d195804;
#10 word0='d195841;
#10 word0='d195878;
#10 word0='d195915;
#10 word0='d195952;
#10 word0='d195989;
#10 word0='d196026;
#10 word0='d196063;
#10 word0='d196100;
#10 word0='d196137;
#10 word0='d196174;
#10 word0='d196211;
#10 word0='d196248;
#10 word0='d196285;
#10 word0='d196322;
#10 word0='d196359;
#10 word0='d196396;
#10 word0='d196433;
#10 word0='d196470;
#10 word0='d196507;
#10 word0='d196544;
#10 word0='d196581;
#10 word0='d196618;
#10 word0='d196655;
#10 word0='d196692;
#10 word0='d196729;
#10 word0='d196766;
#10 word0='d196803;
#10 word0='d196840;
#10 word0='d196877;
#10 word0='d196914;
#10 word0='d196951;
#10 word0='d196988;
#10 word0='d197025;
#10 word0='d197062;
#10 word0='d197099;
#10 word0='d197136;
#10 word0='d197173;
#10 word0='d197210;
#10 word0='d197247;
#10 word0='d197284;
#10 word0='d197321;
#10 word0='d197358;
#10 word0='d197395;
#10 word0='d197432;
#10 word0='d197469;
#10 word0='d197506;
#10 word0='d197543;
#10 word0='d197580;
#10 word0='d197617;
#10 word0='d197654;
#10 word0='d197691;
#10 word0='d197728;
#10 word0='d197765;
#10 word0='d197802;
#10 word0='d197839;
#10 word0='d197876;
#10 word0='d197913;
#10 word0='d197950;
#10 word0='d197987;
#10 word0='d198024;
#10 word0='d198061;
#10 word0='d198098;
#10 word0='d198135;
#10 word0='d198172;
#10 word0='d198209;
#10 word0='d198246;
#10 word0='d198283;
#10 word0='d198320;
#10 word0='d198357;
#10 word0='d198394;
#10 word0='d198431;
#10 word0='d198468;
#10 word0='d198505;
#10 word0='d198542;
#10 word0='d198579;
#10 word0='d198616;
#10 word0='d198653;
#10 word0='d198690;
#10 word0='d198727;
#10 word0='d198764;
#10 word0='d198801;
#10 word0='d198838;
#10 word0='d198875;
#10 word0='d198912;
#10 word0='d198949;
#10 word0='d198986;
#10 word0='d199023;
#10 word0='d199060;
#10 word0='d199097;
#10 word0='d199134;
#10 word0='d199171;
#10 word0='d199208;
#10 word0='d199245;
#10 word0='d199282;
#10 word0='d199319;
#10 word0='d199356;
#10 word0='d199393;
#10 word0='d199430;
#10 word0='d199467;
#10 word0='d199504;
#10 word0='d199541;
#10 word0='d199578;
#10 word0='d199615;
#10 word0='d199652;
#10 word0='d199689;
#10 word0='d199726;
#10 word0='d199763;
#10 word0='d199800;
#10 word0='d199837;
#10 word0='d199874;
#10 word0='d199911;
#10 word0='d199948;
#10 word0='d199985;
#10 word0='d200022;
#10 word0='d200059;
#10 word0='d200096;
#10 word0='d200133;
#10 word0='d200170;
#10 word0='d200207;
#10 word0='d200244;
#10 word0='d200281;
#10 word0='d200318;
#10 word0='d200355;
#10 word0='d200392;
#10 word0='d200429;
#10 word0='d200466;
#10 word0='d200503;
#10 word0='d200540;
#10 word0='d200577;
#10 word0='d200614;
#10 word0='d200651;
#10 word0='d200688;
#10 word0='d200725;
#10 word0='d200762;
#10 word0='d200799;
#10 word0='d200836;
#10 word0='d200873;
#10 word0='d200910;
#10 word0='d200947;
#10 word0='d200984;
#10 word0='d201021;
#10 word0='d201058;
#10 word0='d201095;
#10 word0='d201132;
#10 word0='d201169;
#10 word0='d201206;
#10 word0='d201243;
#10 word0='d201280;
#10 word0='d201317;
#10 word0='d201354;
#10 word0='d201391;
#10 word0='d201428;
#10 word0='d201465;
#10 word0='d201502;
#10 word0='d201539;
#10 word0='d201576;
#10 word0='d201613;
#10 word0='d201650;
#10 word0='d201687;
#10 word0='d201724;
#10 word0='d201761;
#10 word0='d201798;
#10 word0='d201835;
#10 word0='d201872;
#10 word0='d201909;
#10 word0='d201946;
#10 word0='d201983;
#10 word0='d202020;
#10 word0='d202057;
#10 word0='d202094;
#10 word0='d202131;
#10 word0='d202168;
#10 word0='d202205;
#10 word0='d202242;
#10 word0='d202279;
#10 word0='d202316;
#10 word0='d202353;
#10 word0='d202390;
#10 word0='d202427;
#10 word0='d202464;
#10 word0='d202501;
#10 word0='d202538;
#10 word0='d202575;
#10 word0='d202612;
#10 word0='d202649;
#10 word0='d202686;
#10 word0='d202723;
#10 word0='d202760;
#10 word0='d202797;
#10 word0='d202834;
#10 word0='d202871;
#10 word0='d202908;
#10 word0='d202945;
#10 word0='d202982;
#10 word0='d203019;
#10 word0='d203056;
#10 word0='d203093;
#10 word0='d203130;
#10 word0='d203167;
#10 word0='d203204;
#10 word0='d203241;
#10 word0='d203278;
#10 word0='d203315;
#10 word0='d203352;
#10 word0='d203389;
#10 word0='d203426;
#10 word0='d203463;
#10 word0='d203500;
#10 word0='d203537;
#10 word0='d203574;
#10 word0='d203611;
#10 word0='d203648;
#10 word0='d203685;
#10 word0='d203722;
#10 word0='d203759;
#10 word0='d203796;
#10 word0='d203833;
#10 word0='d203870;
#10 word0='d203907;
#10 word0='d203944;
#10 word0='d203981;
#10 word0='d204018;
#10 word0='d204055;
#10 word0='d204092;
#10 word0='d204129;
#10 word0='d204166;
#10 word0='d204203;
#10 word0='d204240;
#10 word0='d204277;
#10 word0='d204314;
#10 word0='d204351;
#10 word0='d204388;
#10 word0='d204425;
#10 word0='d204462;
#10 word0='d204499;
#10 word0='d204536;
#10 word0='d204573;
#10 word0='d204610;
#10 word0='d204647;
#10 word0='d204684;
#10 word0='d204721;
#10 word0='d204758;
#10 word0='d204795;
#10 word0='d204832;
#10 word0='d204869;
#10 word0='d204906;
#10 word0='d204943;
#10 word0='d204980;
#10 word0='d205017;
#10 word0='d205054;
#10 word0='d205091;
#10 word0='d205128;
#10 word0='d205165;
#10 word0='d205202;
#10 word0='d205239;
#10 word0='d205276;
#10 word0='d205313;
#10 word0='d205350;
#10 word0='d205387;
#10 word0='d205424;
#10 word0='d205461;
#10 word0='d205498;
#10 word0='d205535;
#10 word0='d205572;
#10 word0='d205609;
#10 word0='d205646;
#10 word0='d205683;
#10 word0='d205720;
#10 word0='d205757;
#10 word0='d205794;
#10 word0='d205831;
#10 word0='d205868;
#10 word0='d205905;
#10 word0='d205942;
#10 word0='d205979;
#10 word0='d206016;
#10 word0='d206053;
#10 word0='d206090;
#10 word0='d206127;
#10 word0='d206164;
#10 word0='d206201;
#10 word0='d206238;
#10 word0='d206275;
#10 word0='d206312;
#10 word0='d206349;
#10 word0='d206386;
#10 word0='d206423;
#10 word0='d206460;
#10 word0='d206497;
#10 word0='d206534;
#10 word0='d206571;
#10 word0='d206608;
#10 word0='d206645;
#10 word0='d206682;
#10 word0='d206719;
#10 word0='d206756;
#10 word0='d206793;
#10 word0='d206830;
#10 word0='d206867;
#10 word0='d206904;
#10 word0='d206941;
#10 word0='d206978;
#10 word0='d207015;
#10 word0='d207052;
#10 word0='d207089;
#10 word0='d207126;
#10 word0='d207163;
#10 word0='d207200;
#10 word0='d207237;
#10 word0='d207274;
#10 word0='d207311;
#10 word0='d207348;
#10 word0='d207385;
#10 word0='d207422;
#10 word0='d207459;
#10 word0='d207496;
#10 word0='d207533;
#10 word0='d207570;
#10 word0='d207607;
#10 word0='d207644;
#10 word0='d207681;
#10 word0='d207718;
#10 word0='d207755;
#10 word0='d207792;
#10 word0='d207829;
#10 word0='d207866;
#10 word0='d207903;
#10 word0='d207940;
#10 word0='d207977;
#10 word0='d208014;
#10 word0='d208051;
#10 word0='d208088;
#10 word0='d208125;
#10 word0='d208162;
#10 word0='d208199;
#10 word0='d208236;
#10 word0='d208273;
#10 word0='d208310;
#10 word0='d208347;
#10 word0='d208384;
#10 word0='d208421;
#10 word0='d208458;
#10 word0='d208495;
#10 word0='d208532;
#10 word0='d208569;
#10 word0='d208606;
#10 word0='d208643;
#10 word0='d208680;
#10 word0='d208717;
#10 word0='d208754;
#10 word0='d208791;
#10 word0='d208828;
#10 word0='d208865;
#10 word0='d208902;
#10 word0='d208939;
#10 word0='d208976;
#10 word0='d209013;
#10 word0='d209050;
#10 word0='d209087;
#10 word0='d209124;
#10 word0='d209161;
#10 word0='d209198;
#10 word0='d209235;
#10 word0='d209272;
#10 word0='d209309;
#10 word0='d209346;
#10 word0='d209383;
#10 word0='d209420;
#10 word0='d209457;
#10 word0='d209494;
#10 word0='d209531;
#10 word0='d209568;
#10 word0='d209605;
#10 word0='d209642;
#10 word0='d209679;
#10 word0='d209716;
#10 word0='d209753;
#10 word0='d209790;
#10 word0='d209827;
#10 word0='d209864;
#10 word0='d209901;
#10 word0='d209938;
#10 word0='d209975;
#10 word0='d210012;
#10 word0='d210049;
#10 word0='d210086;
#10 word0='d210123;
#10 word0='d210160;
#10 word0='d210197;
#10 word0='d210234;
#10 word0='d210271;
#10 word0='d210308;
#10 word0='d210345;
#10 word0='d210382;
#10 word0='d210419;
#10 word0='d210456;
#10 word0='d210493;
#10 word0='d210530;
#10 word0='d210567;
#10 word0='d210604;
#10 word0='d210641;
#10 word0='d210678;
#10 word0='d210715;
#10 word0='d210752;
#10 word0='d210789;
#10 word0='d210826;
#10 word0='d210863;
#10 word0='d210900;
#10 word0='d210937;
#10 word0='d210974;
#10 word0='d211011;
#10 word0='d211048;
#10 word0='d211085;
#10 word0='d211122;
#10 word0='d211159;
#10 word0='d211196;
#10 word0='d211233;
#10 word0='d211270;
#10 word0='d211307;
#10 word0='d211344;
#10 word0='d211381;
#10 word0='d211418;
#10 word0='d211455;
#10 word0='d211492;
#10 word0='d211529;
#10 word0='d211566;
#10 word0='d211603;
#10 word0='d211640;
#10 word0='d211677;
#10 word0='d211714;
#10 word0='d211751;
#10 word0='d211788;
#10 word0='d211825;
#10 word0='d211862;
#10 word0='d211899;
#10 word0='d211936;
#10 word0='d211973;
#10 word0='d212010;
#10 word0='d212047;
#10 word0='d212084;
#10 word0='d212121;
#10 word0='d212158;
#10 word0='d212195;
#10 word0='d212232;
#10 word0='d212269;
#10 word0='d212306;
#10 word0='d212343;
#10 word0='d212380;
#10 word0='d212417;
#10 word0='d212454;
#10 word0='d212491;
#10 word0='d212528;
#10 word0='d212565;
#10 word0='d212602;
#10 word0='d212639;
#10 word0='d212676;
#10 word0='d212713;
#10 word0='d212750;
#10 word0='d212787;
#10 word0='d212824;
#10 word0='d212861;
#10 word0='d212898;
#10 word0='d212935;
#10 word0='d212972;
#10 word0='d213009;
#10 word0='d213046;
#10 word0='d213083;
#10 word0='d213120;
#10 word0='d213157;
#10 word0='d213194;
#10 word0='d213231;
#10 word0='d213268;
#10 word0='d213305;
#10 word0='d213342;
#10 word0='d213379;
#10 word0='d213416;
#10 word0='d213453;
#10 word0='d213490;
#10 word0='d213527;
#10 word0='d213564;
#10 word0='d213601;
#10 word0='d213638;
#10 word0='d213675;
#10 word0='d213712;
#10 word0='d213749;
#10 word0='d213786;
#10 word0='d213823;
#10 word0='d213860;
#10 word0='d213897;
#10 word0='d213934;
#10 word0='d213971;
#10 word0='d214008;
#10 word0='d214045;
#10 word0='d214082;
#10 word0='d214119;
#10 word0='d214156;
#10 word0='d214193;
#10 word0='d214230;
#10 word0='d214267;
#10 word0='d214304;
#10 word0='d214341;
#10 word0='d214378;
#10 word0='d214415;
#10 word0='d214452;
#10 word0='d214489;
#10 word0='d214526;
#10 word0='d214563;
#10 word0='d214600;
#10 word0='d214637;
#10 word0='d214674;
#10 word0='d214711;
#10 word0='d214748;
#10 word0='d214785;
#10 word0='d214822;
#10 word0='d214859;
#10 word0='d214896;
#10 word0='d214933;
#10 word0='d214970;
#10 word0='d215007;
#10 word0='d215044;
#10 word0='d215081;
#10 word0='d215118;
#10 word0='d215155;
#10 word0='d215192;
#10 word0='d215229;
#10 word0='d215266;
#10 word0='d215303;
#10 word0='d215340;
#10 word0='d215377;
#10 word0='d215414;
#10 word0='d215451;
#10 word0='d215488;
#10 word0='d215525;
#10 word0='d215562;
#10 word0='d215599;
#10 word0='d215636;
#10 word0='d215673;
#10 word0='d215710;
#10 word0='d215747;
#10 word0='d215784;
#10 word0='d215821;
#10 word0='d215858;
#10 word0='d215895;
#10 word0='d215932;
#10 word0='d215969;
#10 word0='d216006;
#10 word0='d216043;
#10 word0='d216080;
#10 word0='d216117;
#10 word0='d216154;
#10 word0='d216191;
#10 word0='d216228;
#10 word0='d216265;
#10 word0='d216302;
#10 word0='d216339;
#10 word0='d216376;
#10 word0='d216413;
#10 word0='d216450;
#10 word0='d216487;
#10 word0='d216524;
#10 word0='d216561;
#10 word0='d216598;
#10 word0='d216635;
#10 word0='d216672;
#10 word0='d216709;
#10 word0='d216746;
#10 word0='d216783;
#10 word0='d216820;
#10 word0='d216857;
#10 word0='d216894;
#10 word0='d216931;
#10 word0='d216968;
#10 word0='d217005;
#10 word0='d217042;
#10 word0='d217079;
#10 word0='d217116;
#10 word0='d217153;
#10 word0='d217190;
#10 word0='d217227;
#10 word0='d217264;
#10 word0='d217301;
#10 word0='d217338;
#10 word0='d217375;
#10 word0='d217412;
#10 word0='d217449;
#10 word0='d217486;
#10 word0='d217523;
#10 word0='d217560;
#10 word0='d217597;
#10 word0='d217634;
#10 word0='d217671;
#10 word0='d217708;
#10 word0='d217745;
#10 word0='d217782;
#10 word0='d217819;
#10 word0='d217856;
#10 word0='d217893;
#10 word0='d217930;
#10 word0='d217967;
#10 word0='d218004;
#10 word0='d218041;
#10 word0='d218078;
#10 word0='d218115;
#10 word0='d218152;
#10 word0='d218189;
#10 word0='d218226;
#10 word0='d218263;
#10 word0='d218300;
#10 word0='d218337;
#10 word0='d218374;
#10 word0='d218411;
#10 word0='d218448;
#10 word0='d218485;
#10 word0='d218522;
#10 word0='d218559;
#10 word0='d218596;
#10 word0='d218633;
#10 word0='d218670;
#10 word0='d218707;
#10 word0='d218744;
#10 word0='d218781;
#10 word0='d218818;
#10 word0='d218855;
#10 word0='d218892;
#10 word0='d218929;
#10 word0='d218966;
#10 word0='d219003;
#10 word0='d219040;
#10 word0='d219077;
#10 word0='d219114;
#10 word0='d219151;
#10 word0='d219188;
#10 word0='d219225;
#10 word0='d219262;
#10 word0='d219299;
#10 word0='d219336;
#10 word0='d219373;
#10 word0='d219410;
#10 word0='d219447;
#10 word0='d219484;
#10 word0='d219521;
#10 word0='d219558;
#10 word0='d219595;
#10 word0='d219632;
#10 word0='d219669;
#10 word0='d219706;
#10 word0='d219743;
#10 word0='d219780;
#10 word0='d219817;
#10 word0='d219854;
#10 word0='d219891;
#10 word0='d219928;
#10 word0='d219965;
#10 word0='d220002;
#10 word0='d220039;
#10 word0='d220076;
#10 word0='d220113;
#10 word0='d220150;
#10 word0='d220187;
#10 word0='d220224;
#10 word0='d220261;
#10 word0='d220298;
#10 word0='d220335;
#10 word0='d220372;
#10 word0='d220409;
#10 word0='d220446;
#10 word0='d220483;
#10 word0='d220520;
#10 word0='d220557;
#10 word0='d220594;
#10 word0='d220631;
#10 word0='d220668;
#10 word0='d220705;
#10 word0='d220742;
#10 word0='d220779;
#10 word0='d220816;
#10 word0='d220853;
#10 word0='d220890;
#10 word0='d220927;
#10 word0='d220964;
#10 word0='d221001;
#10 word0='d221038;
#10 word0='d221075;
#10 word0='d221112;
#10 word0='d221149;
#10 word0='d221186;
#10 word0='d221223;
#10 word0='d221260;
#10 word0='d221297;
#10 word0='d221334;
#10 word0='d221371;
#10 word0='d221408;
#10 word0='d221445;
#10 word0='d221482;
#10 word0='d221519;
#10 word0='d221556;
#10 word0='d221593;
#10 word0='d221630;
#10 word0='d221667;
#10 word0='d221704;
#10 word0='d221741;
#10 word0='d221778;
#10 word0='d221815;
#10 word0='d221852;
#10 word0='d221889;
#10 word0='d221926;
#10 word0='d221963;
#10 word0='d222000;
#10 word0='d222037;
#10 word0='d222074;
#10 word0='d222111;
#10 word0='d222148;
#10 word0='d222185;
#10 word0='d222222;
#10 word0='d222259;
#10 word0='d222296;
#10 word0='d222333;
#10 word0='d222370;
#10 word0='d222407;
#10 word0='d222444;
#10 word0='d222481;
#10 word0='d222518;
#10 word0='d222555;
#10 word0='d222592;
#10 word0='d222629;
#10 word0='d222666;
#10 word0='d222703;
#10 word0='d222740;
#10 word0='d222777;
#10 word0='d222814;
#10 word0='d222851;
#10 word0='d222888;
#10 word0='d222925;
#10 word0='d222962;
#10 word0='d222999;
#10 word0='d223036;
#10 word0='d223073;
#10 word0='d223110;
#10 word0='d223147;
#10 word0='d223184;
#10 word0='d223221;
#10 word0='d223258;
#10 word0='d223295;
#10 word0='d223332;
#10 word0='d223369;
#10 word0='d223406;
#10 word0='d223443;
#10 word0='d223480;
#10 word0='d223517;
#10 word0='d223554;
#10 word0='d223591;
#10 word0='d223628;
#10 word0='d223665;
#10 word0='d223702;
#10 word0='d223739;
#10 word0='d223776;
#10 word0='d223813;
#10 word0='d223850;
#10 word0='d223887;
#10 word0='d223924;
#10 word0='d223961;
#10 word0='d223998;
#10 word0='d224035;
#10 word0='d224072;
#10 word0='d224109;
#10 word0='d224146;
#10 word0='d224183;
#10 word0='d224220;
#10 word0='d224257;
#10 word0='d224294;
#10 word0='d224331;
#10 word0='d224368;
#10 word0='d224405;
#10 word0='d224442;
#10 word0='d224479;
#10 word0='d224516;
#10 word0='d224553;
#10 word0='d224590;
#10 word0='d224627;
#10 word0='d224664;
#10 word0='d224701;
#10 word0='d224738;
#10 word0='d224775;
#10 word0='d224812;
#10 word0='d224849;
#10 word0='d224886;
#10 word0='d224923;
#10 word0='d224960;
#10 word0='d224997;
#10 word0='d225034;
#10 word0='d225071;
#10 word0='d225108;
#10 word0='d225145;
#10 word0='d225182;
#10 word0='d225219;
#10 word0='d225256;
#10 word0='d225293;
#10 word0='d225330;
#10 word0='d225367;
#10 word0='d225404;
#10 word0='d225441;
#10 word0='d225478;
#10 word0='d225515;
#10 word0='d225552;
#10 word0='d225589;
#10 word0='d225626;
#10 word0='d225663;
#10 word0='d225700;
#10 word0='d225737;
#10 word0='d225774;
#10 word0='d225811;
#10 word0='d225848;
#10 word0='d225885;
#10 word0='d225922;
#10 word0='d225959;
#10 word0='d225996;
#10 word0='d226033;
#10 word0='d226070;
#10 word0='d226107;
#10 word0='d226144;
#10 word0='d226181;
#10 word0='d226218;
#10 word0='d226255;
#10 word0='d226292;
#10 word0='d226329;
#10 word0='d226366;
#10 word0='d226403;
#10 word0='d226440;
#10 word0='d226477;
#10 word0='d226514;
#10 word0='d226551;
#10 word0='d226588;
#10 word0='d226625;
#10 word0='d226662;
#10 word0='d226699;
#10 word0='d226736;
#10 word0='d226773;
#10 word0='d226810;
#10 word0='d226847;
#10 word0='d226884;
#10 word0='d226921;
#10 word0='d226958;
#10 word0='d226995;
#10 word0='d227032;
#10 word0='d227069;
#10 word0='d227106;
#10 word0='d227143;
#10 word0='d227180;
#10 word0='d227217;
#10 word0='d227254;
#10 word0='d227291;
#10 word0='d227328;
#10 word0='d227365;
#10 word0='d227402;
#10 word0='d227439;
#10 word0='d227476;
#10 word0='d227513;
#10 word0='d227550;
#10 word0='d227587;
#10 word0='d227624;
#10 word0='d227661;
#10 word0='d227698;
#10 word0='d227735;
#10 word0='d227772;
#10 word0='d227809;
#10 word0='d227846;
#10 word0='d227883;
#10 word0='d227920;
#10 word0='d227957;
#10 word0='d227994;
#10 word0='d228031;
#10 word0='d228068;
#10 word0='d228105;
#10 word0='d228142;
#10 word0='d228179;
#10 word0='d228216;
#10 word0='d228253;
#10 word0='d228290;
#10 word0='d228327;
#10 word0='d228364;
#10 word0='d228401;
#10 word0='d228438;
#10 word0='d228475;
#10 word0='d228512;
#10 word0='d228549;
#10 word0='d228586;
#10 word0='d228623;
#10 word0='d228660;
#10 word0='d228697;
#10 word0='d228734;
#10 word0='d228771;
#10 word0='d228808;
#10 word0='d228845;
#10 word0='d228882;
#10 word0='d228919;
#10 word0='d228956;
#10 word0='d228993;
#10 word0='d229030;
#10 word0='d229067;
#10 word0='d229104;
#10 word0='d229141;
#10 word0='d229178;
#10 word0='d229215;
#10 word0='d229252;
#10 word0='d229289;
#10 word0='d229326;
#10 word0='d229363;
#10 word0='d229400;
#10 word0='d229437;
#10 word0='d229474;
#10 word0='d229511;
#10 word0='d229548;
#10 word0='d229585;
#10 word0='d229622;
#10 word0='d229659;
#10 word0='d229696;
#10 word0='d229733;
#10 word0='d229770;
#10 word0='d229807;
#10 word0='d229844;
#10 word0='d229881;
#10 word0='d229918;
#10 word0='d229955;
#10 word0='d229992;
#10 word0='d230029;
#10 word0='d230066;
#10 word0='d230103;
#10 word0='d230140;
#10 word0='d230177;
#10 word0='d230214;
#10 word0='d230251;
#10 word0='d230288;
#10 word0='d230325;
#10 word0='d230362;
#10 word0='d230399;
#10 word0='d230436;
#10 word0='d230473;
#10 word0='d230510;
#10 word0='d230547;
#10 word0='d230584;
#10 word0='d230621;
#10 word0='d230658;
#10 word0='d230695;
#10 word0='d230732;
#10 word0='d230769;
#10 word0='d230806;
#10 word0='d230843;
#10 word0='d230880;
#10 word0='d230917;
#10 word0='d230954;
#10 word0='d230991;
#10 word0='d231028;
#10 word0='d231065;
#10 word0='d231102;
#10 word0='d231139;
#10 word0='d231176;
#10 word0='d231213;
#10 word0='d231250;
#10 word0='d231287;
#10 word0='d231324;
#10 word0='d231361;
#10 word0='d231398;
#10 word0='d231435;
#10 word0='d231472;
#10 word0='d231509;
#10 word0='d231546;
#10 word0='d231583;
#10 word0='d231620;
#10 word0='d231657;
#10 word0='d231694;
#10 word0='d231731;
#10 word0='d231768;
#10 word0='d231805;
#10 word0='d231842;
#10 word0='d231879;
#10 word0='d231916;
#10 word0='d231953;
#10 word0='d231990;
#10 word0='d232027;
#10 word0='d232064;
#10 word0='d232101;
#10 word0='d232138;
#10 word0='d232175;
#10 word0='d232212;
#10 word0='d232249;
#10 word0='d232286;
#10 word0='d232323;
#10 word0='d232360;
#10 word0='d232397;
#10 word0='d232434;
#10 word0='d232471;
#10 word0='d232508;
#10 word0='d232545;
#10 word0='d232582;
#10 word0='d232619;
#10 word0='d232656;
#10 word0='d232693;
#10 word0='d232730;
#10 word0='d232767;
#10 word0='d232804;
#10 word0='d232841;
#10 word0='d232878;
#10 word0='d232915;
#10 word0='d232952;
#10 word0='d232989;
#10 word0='d233026;
#10 word0='d233063;
#10 word0='d233100;
#10 word0='d233137;
#10 word0='d233174;
#10 word0='d233211;
#10 word0='d233248;
#10 word0='d233285;
#10 word0='d233322;
#10 word0='d233359;
#10 word0='d233396;
#10 word0='d233433;
#10 word0='d233470;
#10 word0='d233507;
#10 word0='d233544;
#10 word0='d233581;
#10 word0='d233618;
#10 word0='d233655;
#10 word0='d233692;
#10 word0='d233729;
#10 word0='d233766;
#10 word0='d233803;
#10 word0='d233840;
#10 word0='d233877;
#10 word0='d233914;
#10 word0='d233951;
#10 word0='d233988;
#10 word0='d234025;
#10 word0='d234062;
#10 word0='d234099;
#10 word0='d234136;
#10 word0='d234173;
#10 word0='d234210;
#10 word0='d234247;
#10 word0='d234284;
#10 word0='d234321;
#10 word0='d234358;
#10 word0='d234395;
#10 word0='d234432;
#10 word0='d234469;
#10 word0='d234506;
#10 word0='d234543;
#10 word0='d234580;
#10 word0='d234617;
#10 word0='d234654;
#10 word0='d234691;
#10 word0='d234728;
#10 word0='d234765;
#10 word0='d234802;
#10 word0='d234839;
#10 word0='d234876;
#10 word0='d234913;
#10 word0='d234950;
#10 word0='d234987;
#10 word0='d235024;
#10 word0='d235061;
#10 word0='d235098;
#10 word0='d235135;
#10 word0='d235172;
#10 word0='d235209;
#10 word0='d235246;
#10 word0='d235283;
#10 word0='d235320;
#10 word0='d235357;
#10 word0='d235394;
#10 word0='d235431;
#10 word0='d235468;
#10 word0='d235505;
#10 word0='d235542;
#10 word0='d235579;
#10 word0='d235616;
#10 word0='d235653;
#10 word0='d235690;
#10 word0='d235727;
#10 word0='d235764;
#10 word0='d235801;
#10 word0='d235838;
#10 word0='d235875;
#10 word0='d235912;
#10 word0='d235949;
#10 word0='d235986;
#10 word0='d236023;
#10 word0='d236060;
#10 word0='d236097;
#10 word0='d236134;
#10 word0='d236171;
#10 word0='d236208;
#10 word0='d236245;
#10 word0='d236282;
#10 word0='d236319;
#10 word0='d236356;
#10 word0='d236393;
#10 word0='d236430;
#10 word0='d236467;
#10 word0='d236504;
#10 word0='d236541;
#10 word0='d236578;
#10 word0='d236615;
#10 word0='d236652;
#10 word0='d236689;
#10 word0='d236726;
#10 word0='d236763;
#10 word0='d236800;
#10 word0='d236837;
#10 word0='d236874;
#10 word0='d236911;
#10 word0='d236948;
#10 word0='d236985;
#10 word0='d237022;
#10 word0='d237059;
#10 word0='d237096;
#10 word0='d237133;
#10 word0='d237170;
#10 word0='d237207;
#10 word0='d237244;
#10 word0='d237281;
#10 word0='d237318;
#10 word0='d237355;
#10 word0='d237392;
#10 word0='d237429;
#10 word0='d237466;
#10 word0='d237503;
#10 word0='d237540;
#10 word0='d237577;
#10 word0='d237614;
#10 word0='d237651;
#10 word0='d237688;
#10 word0='d237725;
#10 word0='d237762;
#10 word0='d237799;
#10 word0='d237836;
#10 word0='d237873;
#10 word0='d237910;
#10 word0='d237947;
#10 word0='d237984;
#10 word0='d238021;
#10 word0='d238058;
#10 word0='d238095;
#10 word0='d238132;
#10 word0='d238169;
#10 word0='d238206;
#10 word0='d238243;
#10 word0='d238280;
#10 word0='d238317;
#10 word0='d238354;
#10 word0='d238391;
#10 word0='d238428;
#10 word0='d238465;
#10 word0='d238502;
#10 word0='d238539;
#10 word0='d238576;
#10 word0='d238613;
#10 word0='d238650;
#10 word0='d238687;
#10 word0='d238724;
#10 word0='d238761;
#10 word0='d238798;
#10 word0='d238835;
#10 word0='d238872;
#10 word0='d238909;
#10 word0='d238946;
#10 word0='d238983;
#10 word0='d239020;
#10 word0='d239057;
#10 word0='d239094;
#10 word0='d239131;
#10 word0='d239168;
#10 word0='d239205;
#10 word0='d239242;
#10 word0='d239279;
#10 word0='d239316;
#10 word0='d239353;
#10 word0='d239390;
#10 word0='d239427;
#10 word0='d239464;
#10 word0='d239501;
#10 word0='d239538;
#10 word0='d239575;
#10 word0='d239612;
#10 word0='d239649;
#10 word0='d239686;
#10 word0='d239723;
#10 word0='d239760;
#10 word0='d239797;
#10 word0='d239834;
#10 word0='d239871;
#10 word0='d239908;
#10 word0='d239945;
#10 word0='d239982;
#10 word0='d240019;
#10 word0='d240056;
#10 word0='d240093;
#10 word0='d240130;
#10 word0='d240167;
#10 word0='d240204;
#10 word0='d240241;
#10 word0='d240278;
#10 word0='d240315;
#10 word0='d240352;
#10 word0='d240389;
#10 word0='d240426;
#10 word0='d240463;
#10 word0='d240500;
#10 word0='d240537;
#10 word0='d240574;
#10 word0='d240611;
#10 word0='d240648;
#10 word0='d240685;
#10 word0='d240722;
#10 word0='d240759;
#10 word0='d240796;
#10 word0='d240833;
#10 word0='d240870;
#10 word0='d240907;
#10 word0='d240944;
#10 word0='d240981;
#10 word0='d241018;
#10 word0='d241055;
#10 word0='d241092;
#10 word0='d241129;
#10 word0='d241166;
#10 word0='d241203;
#10 word0='d241240;
#10 word0='d241277;
#10 word0='d241314;
#10 word0='d241351;
#10 word0='d241388;
#10 word0='d241425;
#10 word0='d241462;
#10 word0='d241499;
#10 word0='d241536;
#10 word0='d241573;
#10 word0='d241610;
#10 word0='d241647;
#10 word0='d241684;
#10 word0='d241721;
#10 word0='d241758;
#10 word0='d241795;
#10 word0='d241832;
#10 word0='d241869;
#10 word0='d241906;
#10 word0='d241943;
#10 word0='d241980;
#10 word0='d242017;
#10 word0='d242054;
#10 word0='d242091;
#10 word0='d242128;
#10 word0='d242165;
#10 word0='d242202;
#10 word0='d242239;
#10 word0='d242276;
#10 word0='d242313;
#10 word0='d242350;
#10 word0='d242387;
#10 word0='d242424;
#10 word0='d242461;
#10 word0='d242498;
#10 word0='d242535;
#10 word0='d242572;
#10 word0='d242609;
#10 word0='d242646;
#10 word0='d242683;
#10 word0='d242720;
#10 word0='d242757;
#10 word0='d242794;
#10 word0='d242831;
#10 word0='d242868;
#10 word0='d242905;
#10 word0='d242942;
#10 word0='d242979;
#10 word0='d243016;
#10 word0='d243053;
#10 word0='d243090;
#10 word0='d243127;
#10 word0='d243164;
#10 word0='d243201;
#10 word0='d243238;
#10 word0='d243275;
#10 word0='d243312;
#10 word0='d243349;
#10 word0='d243386;
#10 word0='d243423;
#10 word0='d243460;
#10 word0='d243497;
#10 word0='d243534;
#10 word0='d243571;
#10 word0='d243608;
#10 word0='d243645;
#10 word0='d243682;
#10 word0='d243719;
#10 word0='d243756;
#10 word0='d243793;
#10 word0='d243830;
#10 word0='d243867;
#10 word0='d243904;
#10 word0='d243941;
#10 word0='d243978;
#10 word0='d244015;
#10 word0='d244052;
#10 word0='d244089;
#10 word0='d244126;
#10 word0='d244163;
#10 word0='d244200;
#10 word0='d244237;
#10 word0='d244274;
#10 word0='d244311;
#10 word0='d244348;
#10 word0='d244385;
#10 word0='d244422;
#10 word0='d244459;
#10 word0='d244496;
#10 word0='d244533;
#10 word0='d244570;
#10 word0='d244607;
#10 word0='d244644;
#10 word0='d244681;
#10 word0='d244718;
#10 word0='d244755;
#10 word0='d244792;
#10 word0='d244829;
#10 word0='d244866;
#10 word0='d244903;
#10 word0='d244940;
#10 word0='d244977;
#10 word0='d245014;
#10 word0='d245051;
#10 word0='d245088;
#10 word0='d245125;
#10 word0='d245162;
#10 word0='d245199;
#10 word0='d245236;
#10 word0='d245273;
#10 word0='d245310;
#10 word0='d245347;
#10 word0='d245384;
#10 word0='d245421;
#10 word0='d245458;
#10 word0='d245495;
#10 word0='d245532;
#10 word0='d245569;
#10 word0='d245606;
#10 word0='d245643;
#10 word0='d245680;
#10 word0='d245717;
#10 word0='d245754;
#10 word0='d245791;
#10 word0='d245828;
#10 word0='d245865;
#10 word0='d245902;
#10 word0='d245939;
#10 word0='d245976;
#10 word0='d246013;
#10 word0='d246050;
#10 word0='d246087;
#10 word0='d246124;
#10 word0='d246161;
#10 word0='d246198;
#10 word0='d246235;
#10 word0='d246272;
#10 word0='d246309;
#10 word0='d246346;
#10 word0='d246383;
#10 word0='d246420;
#10 word0='d246457;
#10 word0='d246494;
#10 word0='d246531;
#10 word0='d246568;
#10 word0='d246605;
#10 word0='d246642;
#10 word0='d246679;
#10 word0='d246716;
#10 word0='d246753;
#10 word0='d246790;
#10 word0='d246827;
#10 word0='d246864;
#10 word0='d246901;
#10 word0='d246938;
#10 word0='d246975;
#10 word0='d247012;
#10 word0='d247049;
#10 word0='d247086;
#10 word0='d247123;
#10 word0='d247160;
#10 word0='d247197;
#10 word0='d247234;
#10 word0='d247271;
#10 word0='d247308;
#10 word0='d247345;
#10 word0='d247382;
#10 word0='d247419;
#10 word0='d247456;
#10 word0='d247493;
#10 word0='d247530;
#10 word0='d247567;
#10 word0='d247604;
#10 word0='d247641;
#10 word0='d247678;
#10 word0='d247715;
#10 word0='d247752;
#10 word0='d247789;
#10 word0='d247826;
#10 word0='d247863;
#10 word0='d247900;
#10 word0='d247937;
#10 word0='d247974;
#10 word0='d248011;
#10 word0='d248048;
#10 word0='d248085;
#10 word0='d248122;
#10 word0='d248159;
#10 word0='d248196;
#10 word0='d248233;
#10 word0='d248270;
#10 word0='d248307;
#10 word0='d248344;
#10 word0='d248381;
#10 word0='d248418;
#10 word0='d248455;
#10 word0='d248492;
#10 word0='d248529;
#10 word0='d248566;
#10 word0='d248603;
#10 word0='d248640;
#10 word0='d248677;
#10 word0='d248714;
#10 word0='d248751;
#10 word0='d248788;
#10 word0='d248825;
#10 word0='d248862;
#10 word0='d248899;
#10 word0='d248936;
#10 word0='d248973;
#10 word0='d249010;
#10 word0='d249047;
#10 word0='d249084;
#10 word0='d249121;
#10 word0='d249158;
#10 word0='d249195;
#10 word0='d249232;
#10 word0='d249269;
#10 word0='d249306;
#10 word0='d249343;
#10 word0='d249380;
#10 word0='d249417;
#10 word0='d249454;
#10 word0='d249491;
#10 word0='d249528;
#10 word0='d249565;
#10 word0='d249602;
#10 word0='d249639;
#10 word0='d249676;
#10 word0='d249713;
#10 word0='d249750;
#10 word0='d249787;
#10 word0='d249824;
#10 word0='d249861;
#10 word0='d249898;
#10 word0='d249935;
#10 word0='d249972;
#10 word0='d250009;
#10 word0='d250046;
#10 word0='d250083;
#10 word0='d250120;
#10 word0='d250157;
#10 word0='d250194;
#10 word0='d250231;
#10 word0='d250268;
#10 word0='d250305;
#10 word0='d250342;
#10 word0='d250379;
#10 word0='d250416;
#10 word0='d250453;
#10 word0='d250490;
#10 word0='d250527;
#10 word0='d250564;
#10 word0='d250601;
#10 word0='d250638;
#10 word0='d250675;
#10 word0='d250712;
#10 word0='d250749;
#10 word0='d250786;
#10 word0='d250823;
#10 word0='d250860;
#10 word0='d250897;
#10 word0='d250934;
#10 word0='d250971;
#10 word0='d251008;
#10 word0='d251045;
#10 word0='d251082;
#10 word0='d251119;
#10 word0='d251156;
#10 word0='d251193;
#10 word0='d251230;
#10 word0='d251267;
#10 word0='d251304;
#10 word0='d251341;
#10 word0='d251378;
#10 word0='d251415;
#10 word0='d251452;
#10 word0='d251489;
#10 word0='d251526;
#10 word0='d251563;
#10 word0='d251600;
#10 word0='d251637;
#10 word0='d251674;
#10 word0='d251711;
#10 word0='d251748;
#10 word0='d251785;
#10 word0='d251822;
#10 word0='d251859;
#10 word0='d251896;
#10 word0='d251933;
#10 word0='d251970;
#10 word0='d252007;
#10 word0='d252044;
#10 word0='d252081;
#10 word0='d252118;
#10 word0='d252155;
#10 word0='d252192;
#10 word0='d252229;
#10 word0='d252266;
#10 word0='d252303;
#10 word0='d252340;
#10 word0='d252377;
#10 word0='d252414;
#10 word0='d252451;
#10 word0='d252488;
#10 word0='d252525;
#10 word0='d252562;
#10 word0='d252599;
#10 word0='d252636;
#10 word0='d252673;
#10 word0='d252710;
#10 word0='d252747;
#10 word0='d252784;
#10 word0='d252821;
#10 word0='d252858;
#10 word0='d252895;
#10 word0='d252932;
#10 word0='d252969;
#10 word0='d253006;
#10 word0='d253043;
#10 word0='d253080;
#10 word0='d253117;
#10 word0='d253154;
#10 word0='d253191;
#10 word0='d253228;
#10 word0='d253265;
#10 word0='d253302;
#10 word0='d253339;
#10 word0='d253376;
#10 word0='d253413;
#10 word0='d253450;
#10 word0='d253487;
#10 word0='d253524;
#10 word0='d253561;
#10 word0='d253598;
#10 word0='d253635;
#10 word0='d253672;
#10 word0='d253709;
#10 word0='d253746;
#10 word0='d253783;
#10 word0='d253820;
#10 word0='d253857;
#10 word0='d253894;
#10 word0='d253931;
#10 word0='d253968;
#10 word0='d254005;
#10 word0='d254042;
#10 word0='d254079;
#10 word0='d254116;
#10 word0='d254153;
#10 word0='d254190;
#10 word0='d254227;
#10 word0='d254264;
#10 word0='d254301;
#10 word0='d254338;
#10 word0='d254375;
#10 word0='d254412;
#10 word0='d254449;
#10 word0='d254486;
#10 word0='d254523;
#10 word0='d254560;
#10 word0='d254597;
#10 word0='d254634;
#10 word0='d254671;
#10 word0='d254708;
#10 word0='d254745;
#10 word0='d254782;
#10 word0='d254819;
#10 word0='d254856;
#10 word0='d254893;
#10 word0='d254930;
#10 word0='d254967;
#10 word0='d255004;
#10 word0='d255041;
#10 word0='d255078;
#10 word0='d255115;
#10 word0='d255152;
#10 word0='d255189;
#10 word0='d255226;
#10 word0='d255263;
#10 word0='d255300;
#10 word0='d255337;
#10 word0='d255374;
#10 word0='d255411;
#10 word0='d255448;
#10 word0='d255485;
#10 word0='d255522;
#10 word0='d255559;
#10 word0='d255596;
#10 word0='d255633;
#10 word0='d255670;
#10 word0='d255707;
#10 word0='d255744;
#10 word0='d255781;
#10 word0='d255818;
#10 word0='d255855;
#10 word0='d255892;
#10 word0='d255929;
#10 word0='d255966;
#10 word0='d256003;
#10 word0='d256040;
#10 word0='d256077;
#10 word0='d256114;
#10 word0='d256151;
#10 word0='d256188;
#10 word0='d256225;
#10 word0='d256262;
#10 word0='d256299;
#10 word0='d256336;
#10 word0='d256373;
#10 word0='d256410;
#10 word0='d256447;
#10 word0='d256484;
#10 word0='d256521;
#10 word0='d256558;
#10 word0='d256595;
#10 word0='d256632;
#10 word0='d256669;
#10 word0='d256706;
#10 word0='d256743;
#10 word0='d256780;
#10 word0='d256817;
#10 word0='d256854;
#10 word0='d256891;
#10 word0='d256928;
#10 word0='d256965;
#10 word0='d257002;
#10 word0='d257039;
#10 word0='d257076;
#10 word0='d257113;
#10 word0='d257150;
#10 word0='d257187;
#10 word0='d257224;
#10 word0='d257261;
#10 word0='d257298;
#10 word0='d257335;
#10 word0='d257372;
#10 word0='d257409;
#10 word0='d257446;
#10 word0='d257483;
#10 word0='d257520;
#10 word0='d257557;
#10 word0='d257594;
#10 word0='d257631;
#10 word0='d257668;
#10 word0='d257705;
#10 word0='d257742;
#10 word0='d257779;
#10 word0='d257816;
#10 word0='d257853;
#10 word0='d257890;
#10 word0='d257927;
#10 word0='d257964;
#10 word0='d258001;
#10 word0='d258038;
#10 word0='d258075;
#10 word0='d258112;
#10 word0='d258149;
#10 word0='d258186;
#10 word0='d258223;
#10 word0='d258260;
#10 word0='d258297;
#10 word0='d258334;
#10 word0='d258371;
#10 word0='d258408;
#10 word0='d258445;
#10 word0='d258482;
#10 word0='d258519;
#10 word0='d258556;
#10 word0='d258593;
#10 word0='d258630;
#10 word0='d258667;
#10 word0='d258704;
#10 word0='d258741;
#10 word0='d258778;
#10 word0='d258815;
#10 word0='d258852;
#10 word0='d258889;
#10 word0='d258926;
#10 word0='d258963;
#10 word0='d259000;
#10 word0='d259037;
#10 word0='d259074;
#10 word0='d259111;
#10 word0='d259148;
#10 word0='d259185;
#10 word0='d259222;
#10 word0='d259259;
#10 word0='d259296;
#10 word0='d259333;
#10 word0='d259370;
#10 word0='d259407;
#10 word0='d259444;
#10 word0='d259481;
#10 word0='d259518;
#10 word0='d259555;
#10 word0='d259592;
#10 word0='d259629;
#10 word0='d259666;
#10 word0='d259703;
#10 word0='d259740;
#10 word0='d259777;
#10 word0='d259814;
#10 word0='d259851;
#10 word0='d259888;
#10 word0='d259925;
#10 word0='d259962;
#10 word0='d259999;
#10 word0='d260036;
#10 word0='d260073;
#10 word0='d260110;
#10 word0='d260147;
#10 word0='d260184;
#10 word0='d260221;
#10 word0='d260258;
#10 word0='d260295;
#10 word0='d260332;
#10 word0='d260369;
#10 word0='d260406;
#10 word0='d260443;
#10 word0='d260480;
#10 word0='d260517;
#10 word0='d260554;
#10 word0='d260591;
#10 word0='d260628;
#10 word0='d260665;
#10 word0='d260702;
#10 word0='d260739;
#10 word0='d260776;
#10 word0='d260813;
#10 word0='d260850;
#10 word0='d260887;
#10 word0='d260924;
#10 word0='d260961;
#10 word0='d260998;
#10 word0='d261035;
#10 word0='d261072;
#10 word0='d261109;
#10 word0='d261146;
#10 word0='d261183;
#10 word0='d261220;
#10 word0='d261257;
#10 word0='d261294;
#10 word0='d261331;
#10 word0='d261368;
#10 word0='d261405;
#10 word0='d261442;
#10 word0='d261479;
#10 word0='d261516;
#10 word0='d261553;
#10 word0='d261590;
#10 word0='d261627;
#10 word0='d261664;
#10 word0='d261701;
#10 word0='d261738;
#10 word0='d261775;
#10 word0='d261812;
#10 word0='d261849;
#10 word0='d261886;
#10 word0='d261923;
#10 word0='d261960;
#10 word0='d261997;
#10 word0='d262034;
#10 word0='d262071;
#10 word0='d262108;
#20 $stop;
    end   
endmodule
