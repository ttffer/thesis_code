`timescale 1ns/1ps
module tb;
reg clk,rst,valid;
reg [1152-1:0] img;
wire [7:0] number;
top_tcb_144_32_10 top_DUT(
    .clk(clk),
    .rst(rst),
    .img_source(img),
    .valid_top(valid),
    .ready_top(ready_top),
    .number(number)
);
always #5 clk=~clk;
initial 
begin
$monitor("number is %d",number);
clk=0;rst=1'b1;valid=1'b1;
img=1152'b0;
#10 rst=1'b0;
@(negedge clk) #(10/4) img=1152'b001111110101001101010000010000100100100001000001001110100011100000111000001111110100010101001011010010000101000101001001010001100100001100111111001111110100000001000011010101100100010101001011010011110100101001001000010001000011111000111010001110110011111001010100011001000100110101001001010000000100000100111111001101110011001100111111010010100100100001101000010101100101100001010101001000100010011100100110001000000010100100111001010001110011010001000101010001000101011101011010000110110010001000100001001011000010111000101111001100110011100000110001001110100101010101011101000111010010110100101010001101110100000100110010010001000100111000101100001001000100011101010000000110100010011100101001001110010100000000101011001111110100100000111110000111110100010001001011000101100001101100100111001101000011000100100101001100110011110100111111000111100011001101000000000101110001100000100110001100100011011000100011001001000010001100011000000101010001100000100001000101000001011000011110001010010010100100011011000110100010011100011001000101100001011000010110000100010001010000010111000110010001100100010101000101010001100100010110000101110001100000010110001010000011110000111100001011110011010100101111001010010010011100101000001011100010110100110011001100010011100000110010001100000010111100101100001011000010111000110111010010110010111100110010001110010011010000110011001011110010101100101010001010100010110101001100011000110100000100110011001100000011001100101110001010010010100000110100001111110100000001100111010101010101010001001100001101100011011100100110000111110010111000111011010010010011011001000101010000100101011001011010001101100011000100100100001100010011100100110101001110010011111000111011001111010101000101011001001011100011001000101100001110110100011000110111010010000101010100111010001110000100100001001101001000010010100100101100001111010100010000101111010001010100111001000110001110100100101101001000001001010001111100101010001110010011011000100111001101110100010101001110001111010100000001000001001011110010001000101010001101100011101000101000001011110011101000111011001110100011000100101111001100000010111000101000001011100011000100101101001101010100001100111100001110100011100000110111001011110011000100110001001100010011010100111001001110100011100100111001001110100011100100111000000011110010000100100100000110000001111100011011000101000001000100010010000110000001010000011001000110000001101000010111000101100001100000011000000110010001101000100101001111100001100000010100000111110001101100011011000101110001010000010110000110000001101101000001011000010011001100011000000111000001111100011011000110000001101000101001001101110011011101100011010101000101001001000001010000010100000000100100000111010011000000111011010011000011100101000110010000000101010101011010010010000011101100100110001101000100000000111000001111010100010001000001001111100101000001011001001101110011010000101100001111000100100100111001010011000101101101000100010001010100101001001101001001100010100100101101010000000100011000110000010010110101100101010010010011110101000101000110001011110010000100101100001111100011101000101000001111010101000001011101010100010100100001000000010000000010011100101011001110000011110000101010001101100100100101010001010100110100000000111000010000110011110000110000001100010011011100111011010010010101100001010100010100110101001001001100010000000100011001000101010000100100011001010000010101000101001001010000010100010101000101001110;
@(negedge clk) #(10/4) img=1152'b010111110100111101000000001110000010111100100010000100110000101100001001000010000000100100011000010111010100100100111011001011100001111100010110000100000000001000000001000000100000001000010100010101100100001000110101001100000011001000110101001100100000101000000100000011000000100100001010010010010100000000111100001101000010111100110000001100000001110000010011000110100001101100010010010010100100010001000010010001010100101001010001010101000101011001010010010011110100101101000001010101110101011101011000010111010101111101100000011011000111000001101110011000000110000100111011011001100101101001010101010101110110000101100000010101100101001001100110010101100100101100111100011101010110101101100101011010110111001001101001010110100101100101101001011010010110011001011111011110000110111001100101011010110111001101110100011100110111001001110101011100110110010101011101011101110111011101110101011001110110001101101001011100100111010001110110011101100111011001110101011101100111011001110101011011110110101101110010011101010111011001110101011101100111011001110110011101100111010101110101011101010111010101110101011101010111010101110101011101010111010101110110011000010101001101000110001111110011011100100111000110000000111100001101000011100001000100100001010111110100110101000000001100110010000100010010000011000000001000000001000000100000001100011001010110000100001100110101001010110010101000101011001010100000011100000011000010100000100000001100010010000011101000110001001001010001111000011110000111100001000100001011000100100001010100001110010000110011100100110011001101010011100101000000010000010100010001000001001111100011110100110101010100000101000001001111010100110101010101011001011010000110110001101000010110110101110000110001011000110101011001010001010100100101110101011100010100010100110001100011010101000100010100110001011101010110100001100000011010000111000001100110010101100101011001101000011010000110000001011000011110000110110101100010011001110110111001110010011100110111001001110101011100110110001101011001011101110111011101110101011001000101111001100110011100100111001101110110011101100111010101110100011101100111011001110101011011100110100001110010011101010111011001110101011101100111011001110110011101100111010101110101011101010111010001110101011101010111010101110101011101010111010101110110010110100100110101000010001111010011110100110001000111100000110100001100000010110000111100011100010101110100100000111111001110000011010001000001001101000000010000000001000000110000001100010110010100110100001000111010001110100100000101001010010000000000100100000100000011110000100100001011010001100011100100101111001000000001011100010110000101110000111000001001000100000001000100001011001111100011001000101010001011000011000000110111001110010011110000111001001101100011010100101111010010000100011101000110010010100100110001010001011000000110011001100101010110010101011000101110010111000101000001001100010011100101100101011000010010100100010001011110010100010011111100101010011100010110010001011011011000010110101001100001010100000101000001100110011001100101110001010001011101100110100101011100010111110110100001101110011100010111000101110110011100110101110101010000011101110111010101110100010111100101011001100000011100000111001101110111011101100111010001110010011101100111011001110101011011000110010101110000011101010111010101110101011101100111011001110110011101100111010101110101011101000111010001110101011101100111010101110101011101010111010101110110;
@(negedge clk) #(10/4) img=1152'b000010000001011000010111000110000001110100011011000110010001111000011110000110110001100100010111000101000001100100011010000111000010001100100101001001000010001100100010001000000001111000011110000101110001101000100001001001010010101100101111001100110011011000110110001110110100001100111110000110100010001100101100001101110100000000111001010000110100111101000101010010110101010001001101001100010011010101000100010100010101010001001011010100110101101001011000010110010101010001001101010001000100100001010001010011110100111101010110010111000110001001100100010111000100111101001111001011100011101101010010010100010101000001011001010111010101110101011000010010010100001101000100001101010100010001001111010100000100001101000100010011010100101001000101001110100011101000111000010001000100101001000100001110110011111101001000010100110100111101001100010001100100001001000100011010100110100001100001010100000100111001011101011001000110100101101001011001110101101101100010011110000111011101110111011011100110100101110011011100100111000101110010011100010110010001101001011110100111101001111001011101110111100101110111011110010111011101111001011101110110100101101011000010000001001100010011000100110001100000011000000101100001101100011010000110000001010100010100000100010001010100010101000110000001111100100001001000000010000000011110000110110001100100011001000100110001011000011100001000010010011100101010001011010010111100101101001100010011100000110011000101110010000000101000001101000011110000110011001110110100011000111001001111100100011100111111001011100011001101000001010011010101000001000101010010110101000001001011010010110100010000111100010001000100011101001111010011100100101101010000010100110101010101010101010011010100000100111111001011010011101101010011010100010100101001001110010011110101000001001010001111000011100000111000001100100100011101010001010011010011110000111011010000000100000000111101001100110011010000101111010001100100110001000011001101010011011001000000010100000100111101001100010001010011111101000000011011100110110001100010010011010100101001011100011001010110101101101101011010000101100001011111011110000111011101110111011011100110011101110010011100010110111101110001011011010101111001100001011110010111100001111000011101110111011101110101011101100111001001110000011011000101110101011110000001100000111000001101000011110001001000010011000011110001001000010010000100010000111100001110000011010000111100001111000100100001011100011001000101100001011000010101000100100001001000010010000011100000111100010110000110000001111000100000001000110010011000100010001001010010110100100111000100110001100100100000001010110011001100101011001100100011101100101110001100010011100000110000001010110010111100111101010010010100100100111101010000010100001100111110001111100011011000101110010001000100011101001110010011000100011001000110010001010100011101001000010000100011011000110010001010010011110001010110010100100100001101000010010000100100010000111111001100110010111100101100001011010100101001010010010010010011000100101111001101000011011000110110001011000010110000100110010010010100111101000010001011100010110000111000010011010101000101001111010001100011111000111110011100110110111001100010010010000100010001011000011001010110110101110000011010100101011101011011011110010111011101110111011011010110010001110000011100000110111001101110011010000101011101011000011110000111011001110110011101010111010101110010011100110110110101101001011000100101000101010001;
@(negedge clk) #(10/4) img=1152'b001000000010110000100100000111000001111100100000000111110001111100011100000111010001110000011101001010110010001100011101000111000001110000011111000111110001111100011111001000100010010000100011001111010011111001000000001111100011111000111111001111000011100100111011001111110100001000111111011000100110000101010101010011100100111101010111010010000100101001011010011001010110100001100011011010010110010001010001001111010011000000110001001001110010001101000101011011110111000001101011011010110110111001101110011010110110001001011000010000110010111101000110011011100111001001101101011010100110111001101110011011010110110101110000011011100101111001000110010100100110101001101011011010110110111001101110011010110110101001101100011011010110101001100111010111100110010001101001011010110110111001101001010111100101101101011110010111000101101101011100011001010110101001100101011011000110111001100000010101110101010101010101010011110101000101010000010110000110101101100000011010110110111101101001010110000101100001010110010100100101001101010000010111110110110101100001011010000110101101100100011000010110000101011111010111110110000101011101010111010110101001011111001001110011001100101100001000010010001100100101001000110010001000011111000111100001111100100000001100110010100000100000001000000010000000100010001000010010000000100010001000110010001100100101001101110011010000110110001101010011010100110110001101000011010000110110001101110011101000111011010110000101010101001011010001100100011101001111010000010100010001010100010111110110000101011110011000000101110101001101001110010010111000110001001001100010000101000010011010010110101001100111011000100110010001100100011000010101101001010011010000000010111001000011011010010110110001101000011000100110010001100100011001000110010001100111011001000101010101000001010011100110000101100101011001010110011001100100011000010110000101100001011000010101111101011100010101010101101101100001011001000110010101011111010101100101001001010100010100110101001001010010010110010101111001011010011001100110011001011000010011110100110101001100010001110100100101001000010011100101111101010110011001100110011101100000010100010101000001001110010010100100101101001001010101010110000101010111011001010110010101011110010110110101101001011001010110000101101001010101010101010101111001010111001000100010011000100010001000000010010000100101001001000010001100100000001000000001111100100011001001100010000100011111000111110001111100100001001000010010000100100011001001000010010100100111001101000011010000110100001100110011010000110101001100110011001100110101001101110011101000111010010101100101010001001010010001010100011001001111010000100100010001010100010111100110000001011100010111110101110001001100001110010010111000110011001010100010001101000011011010000110100101100110010111100110000001100001010111110101101001010011010000100011000001000011011001110110100101100100010111110110000101100001011000100110001001100101011000110101010001000001010011010101110001100000011000010110001001100000010111100101110001011110010111110101101101011000010100000101010001011100011000000110000101100000010110010101011001011000010101010101001101010101010110010101011001010100011001000110010001100011011000100110001001100001011000000101111001011111011000000101011001001111011001010110011101100100011000100110001101100011011000010110000101011111010111100101100001010000011001000110010101011110010111000101101101011010010110100101101101011000010101010101100101010010;
@(negedge clk) #(10/4) img=1152'b001110110011010000110011001100010010110000110010001111010100011101000001000111110001010000011110001011100010001100100101001111000011111100110001001100010011001101000000001110110001110100100101001011110010101000101111001111110100001100111011001111010011100100110010001111000100001100110111001101110011010000110010001111000100000001001001010001110011010100110010001010110011001100110010001101000010101000110100001111000100001101000111010001010011100000110000001010100010110100110101001000110010111100111101001111000011110100111110001111000011100100111011001101100011001100101101001000000011011100111011001110100011001100110100001100110010110100111000001111010010111100100110000110000011100100111010001011110011000100110011001011110010110100101100001110010011001100100010000110010011110000111100001011010010101100100100000110100010101000011111001010000011001100100001001010000011011101000000001010010001111000011101000111010001110000010011001000100010000100100000001001110010100100110010001001000010001000100011000110100001000100010100001000110010000100101001000111110001100100100111001000100010010100100010000110100001001100010110000111010001011000100001010101010100011101000010001111010011100101001001010111000110010101100000001101100010011000101110010001100011010100110001010001100100100000111111010010100101001101100000010110000011000000110011010001100011110000111011010010000100101101000100010010010100100101001010010110100101101101000110010011010100001101000001010001100100100001010001010100010100001001000001001111100100011000111111010001010011010100111101010001100100101101001110010011000100001000111111001110000011101101000001001100000011101101000101010001110100100001001000010001000100000101000111010001010100000100111010001010110100011001001001010000110011111000111111010000000011100101000101010011000011110000110011001000000100100001001111010000010100001001000100001110110011101100111110010010000100000100101100000111110100100001010010010001110100000000111000001010100011111100101101001100110100000100101110001100110100011101010010001111000010101100101010001100010011000100011100001011000010111100101100001101000011011101000011001100100011001000110011001001110001110000011101001011100011000000110100001010010010011000111000001100000011011100110011001001110001111100011111001010100010000100101011010001010011100100111010001111010011101001000010010010100101010101010001001010100001101000100010001101010010011000110011010100000101001000111100001111000011111101010000010010110010011000101000001011100010111001000011010101010101011001001100010011110011111100111001010010100101000100111100001101000011011101000111010100100101001001011011010110100011110100110010001011110011110000110101001100110010110001000011010100010101011001011010010101100100010000110100001010110010111100110100001001010011010001001100010100010101010001010100010100000100101001000110001101110011001100101110001000110011100001001001010011000100100101001010010010100100001101001000001111100010111100100111000110100011100101000011001111000011111100111110001110110011111000110100001110000011001100100011000110010011101101000100001101100011001000101001001000000011000100100100001010010011001000100000001010100011100001000111001011100010000100011101001000000010000000010100001000010010001100100000001010000010101000111010001001110010010000100101000110110001001000010010000111110010001100101001000111110001110100101110001001010010100100100110000111000001010000010010000110100001100000100010;
@(negedge clk) #(10/4) img=1152'b001001010010001000100111001001010010000100100000001000100010011100101001001010000010101100101001000111110001110000011101000111000001110100100001001001110010010000100110001001110010101100101000001000110001011100001111000010100000110100010011001000000010000100101000001011100010110000101000001001100010101000010011000010110000101000010001000110100001011000010111001011100011000000101011001000000011001100010101000100100001001100100101001010100010111000100010001101110011011100101000000110010010100100010011000101110010111000110101001101000011101100111010001101100011010100100100000110010001101100010101001000010011100000111101001101110011101100110111001101110011001100011111000111010001100000010101000111110010100100101010001101010011100000101011001100010010111100011101000111110001110000011001001000100010010000100101001010110010101000101001001010100010101100101001000111110001101100011001000111000010000000100001001000010010010100101001001010000010101000101110000111000001110000011101000110010001010000011010000111000010000100100101001001000010011100101110000110010001110000010111000101110001010100011010000110100001110100100001001000010010000100100100001010110010100100101110001011010010011100101000001010100010111100110000001011010011000000101111001001000010001100100100001000100010000100100110001011010010101100101110001011100010111100101100001010010001110000010011000011000000111100010111001001010010011100110011001110000011001000101110001011010011001000010111000011010000110100010110000111100001101000011101001101110011011100110000001001010011110000011001000100110001011100101100001100010011011100101000001111110011111100101110000111010011000000010111000111000011011101000000010000000100011101000111010000100011111000101010000111010010001000011001001001100100000101000110010001000100101001000111010001010011111100100110001000100001111100011010001001100011000100110011001111100100100000111110010000110011111000100110001001000010001000100000001100000011000100110010001110000011110000111110001111010011101100110110001001000010000100011111001001110010111000110010001100110011100100111100001110100011110000111101001000010010001000100001000111100001101100101001001011010011001100110111001101010011101000111111000111010010000000011100000111000001101100100100001010010010110100110001001100000011000100110100010010000100011101001110010011010100011101000111010010010101000101001111010011110101001001010010001110110011101000111100001110110011101101000010010011110100100001000111010010110101000001001101001110110010111000011111000100100001100000100111010000100100010001001010010011110101001001010001001110110100010000100111000101010001010100100110001101100010110000101110010010010101000101010010001011110100101100101001001000100010010101000110010011010100101000110110010100000101010101001111001011000100000100100011001010010100100001010101010110010101111001011000010101110101010101001001001100100011010100100101001101000101000101010101010110010101111101011010010111000101011000111011001110100011001100101010001110010100100101000111010011110101101001011000010111010101011100111000001111010011100100110101010010000101001001001111010101010101101101011101010110100101010101001001001111010011101000111001010000100100101101010011010101100101110001011100010110010101010001010001001101110011101000111010001100110010110101000110010100000101011001010111010101000101010001010110001011100011010100101111001011110010110000111001010001010100110101010000010011110100100101001011;
@(negedge clk) #(10/4) img=1152'b000011010000011100000110000100000001010100010001000110000001101100011011001001010010001000010111000010000000011000001010000110000010000100100010001011010010101000011111001000000001111100010000000010010001011100101110000110010010001101000101011000000100010000100101001011010010101000001111000011100011001101001111001001010001110101010010010111000010101000001111001010100011010100010110001011110101000001010111010101010101001101101001010101000001011100010011001001110100000000010011001110000011010000100110010100110111010001101011010001010001101100100010001000010001010000001001000100000001001000100000011001010100111000100011001000010010011000011111000100010000100100000111000001100001000000010011010001000100100000111011001110100010100100010000000001110000011100000110000001010000011100001101000110010010011000011111000110000001000000001000000001100000010100000101000001010000100100001110000110000001000000001000000010000000011100000101000001010000010100000111000001010000100000001100000100010000011100000100000001000000010000000011000000110000011100000111000001000000100100001110000001110000101000000100000000100000001000000010000000100000010000000101000011010000011100000110000011010001001000001111000101010001011100010110001000000001110100010100000010000000010100001001000101000001110100011110001010000010010100011011000111000001101000001110000010100001010000101001000101010001111001000000010110010011110100100000001001110010010000001101000011110010111001000111001000010001100101001100010101010010010100001101001001000010111100010100001011010100101101001111010011110100110101100010010011100001010100010000001000010011110100010100001101000010111100011111010011100110111101100111010000110001101100100000001000000001011000001100000100100001000100011101010111110100101000100010000111110010010000011111000100110000110100001100000010100001001000010100010000100100010100111011001110110010101100010100000011000000101100001010000010110000111000010010000110010010101000100111001000010001100000001110000010110000101000001001000011010001000100010010000110010001100000010011000100010000111000001100000011000000110100010000000010110000110000001110000101110001000100001111000100000001000000010001000100110001101000011110000010100000110100010001000100110001100000010110000110010001101000011111001000100010000100100000000011000000011000000100000010110000111100001100000011110000111000001101000101110001110100100110000010110000010100001000000100110001101100011011001000110001111100010100000101100001111000100110000100110001010000100101000101000001110000111010010100000011010100011010001000000010001100101001000101010010101101000001000111100001011101000110010011000001111000001011000111110010111000111011001100010100011101001101010011000100100001011011010001110001000100001111000111110100101101000111010000000011001000101100010100000110101101100011001111110001101000100000001011000100000101000111001011000001100000011111010110100100011000100011000111110010111000111000010000100100011101000111001101000011000000011011010000010100010101000011010001100100011101000110010001010100011001000101001110010011110000110100000111100100000101010010010100000100110001001000010001100100010101000000001110110011110000101011001000100100000101001000010010100100100101000111010010000100100001001000001110010010110100011110001110000100001101000111010011010101000001010110010111100110010001101010001100110010011100101001010000000100101001010101011000000110010101101111011101010111001001110000;
@(negedge clk) #(10/4) img=1152'b000011010000101100001101000011100000110100001100000100110001100000001111000011110001000100011000000101010001000000010010000110010001010100010000000101010001101000011000000111010010010000100111000101110001010100010100001000010001110100010011000110010001100000100101001100000011010100111100000100010001011100010001000101110001100100010101000110000001010000100000001101110101110001110000000011110001001000001111000101010001110100011011001000000011000100111111010110100111000001101100000101100001100100010001000100000001101100011100001000000011000001000001010011100101001001001000000111100001111100010110000011000001011000011010000101100001101100100011001111000100010101000100001000110010011000011100000011100000111000010010000110000001101100010100001011000100100101001000000111110010001000100001000110000001000000001101000101000001010100001011001000100011100000110000000110100010000000100100001001010010010000010100000010100000101000001101000101110010001100100100000111000001111000011101000111010001111000011010000101100001011100011011001000100010011100101001000100010001001100010100000110010001110100100000001000110010001100100110001010100010100000101010000101110001011100011011000111010001101100011001001000000010010000011010000110010001101000100000001000000001111000101100001101000010110100100111001010000010011000100010001010010010111000101111001000110010010000101111001111110011101100101111001011110010101100110001001101110011101101000010000110100010010100101101001110010011101000110100001100000011010000111000010000110110000001110011000101010010000000110010001110110100000000111110001111010100011001010011011001000111001101110000000111100010101000110011001110000011111000111111001110110011111101010000010101110101100001010000001001010010101100110011001101000011101000111101001110000011000100101110010000110100101101001001001010110011000000110011001101010011010100110111001110110011100100101001001101010100111101001101001010000010101000101110001101110011010100110100001101110011010000101000001011010011111000110110001000000010010100101011001100110011010000110010001100000010110000101001001000000010100100101011000111110010001000100011001001000010010100101000001100010011001000101110001010010010110000101110000100110001010100011000000111010010001000100110001011000011001100110001001011100010110100101111001010010010101100101100001010100010101000101100001011110011001000101011001010100010100100101001001100000010111100101110001011100010101100101001001011000010111100101110001100000011000100110000001100010011010000110010001101010011000000100110001011000010101000110001001101110011100100111110001010110011001000101101001100010011000100101100001011000010101100110000010000000101111001110001001001110010101000101010001100010011010000110011001110100100010001001110011000100111010001110000001011000010111000101011001011010011001000110100001110100100001001010000010101110101100101001110001011000011000100110000001011010011000100110100001100010010110100101111010001000100101001000111001101100011110100110111001011110011000000110000001100000011000000100100001100110100110101001100001101000011010100110100001100110011000000110000001100000010101100011111001010110011110000110011001001100010101000101111001100110011001000110000001010100010010000100000000111100010010100100101001000110010011000100101001001010010010000100101001010110010101100101000001001010010011100101000000100110001010000010101000110100001111100100010001010000010111000101101001010110010100000101001;
@(negedge clk) #(10/4) img=1152'b001110100011011000110110001101100010111100101111001100010100011101011010010010110011111001000011001111010011100000110101001110000011001000111001010000110100110001011010010101100100010101010010001110010011110101000001001111100011101001001010010100100100100001011001010111010100111101011000001101110100000001001000010000000011111101010101010101100101001101100000010111100101010001011100010001010100001001000000001111100100011001001110010111010101110101011011010110100101001101011000010111010101001101000100010000100100011101000001010100110101111001011110010100000100110001010001010111010110011001100111010101100100110101001100010010110101001001010011010010000100111001010011010011100101100101101011010110110100101001000011010001010101010001001110010010110101001101010100010110010101011101101010010111010100100000111001010010000101101001001100010010010100100001000101010111010110000001100011010110010100011100111001001110100100111001010101001111000001110100010100010011000100111101010011010011110011101001000111010000110100010001001110001101110001101000001100010000100100010001000110001111110010101000111101001111000011101000111100001111000010001000001100010000010011110100111101001111010011011000110110001110010100111001100000010101010101001101010101010001000011111100111100001111110011100101000001010011000101000001011111011000010101101101100100010000000100010001000110010001010100001001010001010110010100101101011101011001000110000101101010001111110100011101001110010001110100011101011010010110110101100101100101011001000110000101101100010100000100101001001000010001110100110101010010010111100110000101100001011000000101111001101011011011110110000101010000010010110100111001000111010100110101111101100001010100110101011001100100011011110111010101110110010111110101000101001110010010100101010001011000010100000101101101100101011001000110110101111010011001010100101101000011010001110101010101010010010110000110000101100011011010010110100001110100011001110100101000111010010010100101101001001111010101010101001101010001011010010110101001101011011000100100101100111100001111010100111001010101010010000010000100010110010110100101111001100001010110100011111101010000010011000100101001001111010000110001110100001010010100100101010101010101010010000010111101000111010010110100100101000111010010010010100000001010010010100100011001000110010001100011111001000000010001000101010101100011010101000101000101010011010011010100100001000101010010000100001001001100010101100101110001100100011000000101100001100010010010010100111001001111010011100100101101011011011000100101100101100100011001100101111101100111010010000101000001010111010100000101000001100001011000010110000001101010011010000110000001101010010101110101010001010010010100100101011001011000011000100110001101100100011001010101111101100111011011100110001101010110010100110101010101001110010110000110001001100101011000000101110001100010011010110111001101110110011000010101010001010010010011110101011101011101010111010110000101100101011000010110101001111000011001100100111101001000010011000101100101010111010111010110001101100101011010010110011101110110011010010100111101000000010100000101111101010100010110010101010101010011011011010110110101101111011001000101000001000101010001010101010001011011010100010010010000011000011010100110110001101100010111110100011101011011010101100101000101010110010100100010010000001100011001100110011101101000010101000011011101010100010110110101100101010100010110100011001100001100;
@(negedge clk) #(10/4) img=1152'b011001100011010000100111001111000011010100101010001001100010011100101101010001000101111101100010011000000010110100100010010011000011111100100110000110010010000100110111010001110101110001100100011000000010101100101010010101010100111000100011000110000001101000110100010000110100100001100101011000010011110100111010010001100100000100110001001100010010010100100101001100110011110001100101011001110100010101001011010010000100101001001000001110010011000100101100001100000011111101100011011100010101010101000100001110110100000000111001010000010100000100111101010000010100001001011101011110000110001001001010001110100011111100111111010000110100100001001100010011010100111001100001011110100111011101101000010101010101011001010010010100100101010001000101010100110110100101101111011000110110100001101110011000110110011001100011011000010110000101010101010111000111001101111001010110010101010101100111011000100101110001011111011000100110001101010101011000110111011101111010011000100101110001101010011001010101101101011100010101110101010101010000011000110111100001111001010110010101110101100110011010100110110001101010010111100101100101010110011000100110101101101100010100010010011100011100001011000010011000011110000110110001110100100001001100110100100001001011010011000001111100011001001111000011000100011100000100100001100000101001001101110100100001010000010011100001111000100000010010010100010000011001000100000001001000100111001101000011100001010001010101110010110100101101001101110011001100100101001001000001100100011010001001110011001001011010010111110011001000111000001101010011010100110101001001110010000100011101001001110011011001011101011011000100001000110011001011100011000100101011001011110011000000101010001110100011101101011000011101110101011000111011001010010010100000100110001010000010110000110001010001000100100101011100011110100111011101100100010000110011101100110011001100110011010100101011010000100110010101101100011001100110110001101110010101000100100101000011010000010100010100111010010011010111000101111001011001010110000101101100011000100100011001000000010001000100100100111100010110110111011001111010011011100110101001110001011010110101110101001111010001100100001001000001011000000111100101111001011000100110100001101101011100010111001101101110011000000101100001010111011001000110111101110000010100010010100000011110001011110010100000100000000111010001111000100010001101000100100101001011010011000010000100011011001111100011001100011110000101000001100100101010001110010100101001010010010100000010000000100010010010100100010100011011000100010001001100101000001101110011101001010100010110010010111100101111001110010011010100100111001001010001101100011100001010110011011001011111011000000011010000111010001101100011011100111000001010010010001000011111001010110011101001100011011011010100010000110100001100000011001100101110001100000011001000101100010000010100001001100001011101110101011100111011001010000010100000100110001010000010110000110010010010110101000101100110011110100111011101100100010000010011100000110001001100010011001100101011010001010110100101110001011010010110110101101111010100100100010000111111001111010100001100111001010011100111000101111001011001000110000101101110011000010100001100111100010000000100100000111011010111000111011101111010011010110110100001110001011010110101101001001110010001010100001001000001011000010111100001111001010111110110010101101100011100000111000101101011010111110101101001011001011001100110111101101111;
#100 $finish;
end
endmodule
