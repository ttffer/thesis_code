module layer0_tcbcnn_121_25x64x10
(
    input clk,
    input rst,
    input [475-1:0] layer_in,
    input valid,
    output  reg ready,
    output [27*64-1:0] layer_out
);
parameter DATA_WIDTH = 27;
parameter INPUT_DATA_CNT   =   25;
reg    signed [DATA_WIDTH-1:0]  in_buffer[0:INPUT_DATA_CNT-1];
genvar j;
generate
for(j=0;j<INPUT_DATA_CNT;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=layer_in[j*19+18:j*19+0];
                    end
            end
    end
endgenerate
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0-(0+(in_buffer[0]<<1))-(0+(in_buffer[1]<<4))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<3))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<2))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<3))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<2))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<3))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<2))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<4))-(0+(in_buffer[9]<<2)+(in_buffer[9]<<3))-(0-(in_buffer[10]<<1)+(in_buffer[10]<<4))-(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<5))-(0-(in_buffer[12]<<1)+(in_buffer[12]<<4))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<1))-(0-(in_buffer[14]<<0)+(in_buffer[14]<<3))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<3)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<2)+(in_buffer[17]<<3))-(0-(in_buffer[19]<<0)+(in_buffer[19]<<2)+(in_buffer[19]<<3))-(0+(in_buffer[20]<<1))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<4))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<2))+(0-(in_buffer[23]<<1)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0+(0-(in_buffer[0]<<1)+(in_buffer[0]<<6))-(0+(in_buffer[1]<<5))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<4))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<4))-(0+(in_buffer[4]<<3))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<1)+(in_buffer[5]<<4))+(0+(in_buffer[6]<<1))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<2)+(in_buffer[7]<<6))+(0-(in_buffer[8]<<1)+(in_buffer[8]<<4))+(0-(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<3))+(0-(in_buffer[10]<<0)+(in_buffer[10]<<4))+(0+(in_buffer[11]<<4))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<3)+(in_buffer[12]<<6))+(0-(in_buffer[13]<<2)+(in_buffer[13]<<4)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<6))-(0+(in_buffer[15]<<2)+(in_buffer[15]<<3))-(0+(in_buffer[16]<<1))+(0+(in_buffer[17]<<3)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<4)+(in_buffer[18]<<6))-(0+(in_buffer[19]<<0)-(in_buffer[19]<<2)+(in_buffer[19]<<4)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<4)+(in_buffer[20]<<6))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<5))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<1)+(in_buffer[22]<<6))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<2)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0+(0+(in_buffer[0]<<3))+(0+(in_buffer[1]<<3)+(in_buffer[1]<<4))+(0-(in_buffer[2]<<1)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<1))-(0-(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<3))+(0-(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<4)+(in_buffer[5]<<5))+(0+(in_buffer[6]<<1))-(0+(in_buffer[7]<<1)+(in_buffer[7]<<5))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<3))-(0+(in_buffer[9]<<1)+(in_buffer[9]<<3))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<4))-(0+(in_buffer[11]<<2)+(in_buffer[11]<<5))+(0+(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<6))+(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<4))-(0-(in_buffer[15]<<1)+(in_buffer[15]<<3)+(in_buffer[15]<<4))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<3))+(0+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0-(in_buffer[18]<<1)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<0))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<4))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<4))-(0+(in_buffer[22]<<3)+(in_buffer[22]<<5))-(0-(in_buffer[23]<<0)+(in_buffer[23]<<4))+(0+(in_buffer[24]<<2)+(in_buffer[24]<<4));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<3))-(0-(in_buffer[1]<<0)+(in_buffer[1]<<3)-(in_buffer[1]<<5)+(in_buffer[1]<<8))-(0+(in_buffer[2]<<1)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<4)+(in_buffer[3]<<7))-(0+(in_buffer[4]<<2))+(0+(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<5))-(0+(in_buffer[6]<<1)+(in_buffer[6]<<4)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<1)+(in_buffer[7]<<3)+(in_buffer[7]<<4))+(0-(in_buffer[9]<<1)-(in_buffer[9]<<3)+(in_buffer[9]<<6))-(0+(in_buffer[10]<<4)+(in_buffer[10]<<5))+(0-(in_buffer[11]<<1)+(in_buffer[11]<<4))+(0-(in_buffer[12]<<0)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<3)+(in_buffer[13]<<5))+(0-(in_buffer[14]<<0)+(in_buffer[14]<<5))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<6))+(0+(in_buffer[16]<<0))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<5))+(0+(in_buffer[18]<<2)+(in_buffer[18]<<4)+(in_buffer[18]<<5))-(0+(in_buffer[19]<<2)+(in_buffer[19]<<4)+(in_buffer[19]<<5))+(0-(in_buffer[20]<<0)+(in_buffer[20]<<3))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<3)+(in_buffer[21]<<4))+(0+(in_buffer[22]<<1)-(in_buffer[22]<<3)+(in_buffer[22]<<6))-(0+(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<5))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<4)+(in_buffer[24]<<5)+(in_buffer[24]<<8));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0+(0+(in_buffer[0]<<2)+(in_buffer[0]<<4)+(in_buffer[0]<<5))+(0+(in_buffer[1]<<2))+(0+(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<1)+(in_buffer[3]<<4)+(in_buffer[3]<<6))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<4)+(in_buffer[4]<<6)+(in_buffer[4]<<8))+(0-(in_buffer[5]<<2)+(in_buffer[5]<<4)+(in_buffer[5]<<5))-(0-(in_buffer[6]<<0)-(in_buffer[6]<<2)+(in_buffer[6]<<4)+(in_buffer[6]<<5))+(0+(in_buffer[7]<<1)-(in_buffer[7]<<4)+(in_buffer[7]<<7))-(0+(in_buffer[8]<<3))-(0-(in_buffer[9]<<0)-(in_buffer[9]<<4)+(in_buffer[9]<<9))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<4))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<3)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<1)-(in_buffer[13]<<3)+(in_buffer[13]<<6))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<3))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<3)+(in_buffer[15]<<5))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<3))+(0+(in_buffer[18]<<3))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<2)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<4))+(0+(in_buffer[21]<<3))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<2))-(0+(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0+(0-(in_buffer[0]<<1)-(in_buffer[0]<<4)+(in_buffer[0]<<8))-(0+(in_buffer[1]<<1)+(in_buffer[1]<<3)+(in_buffer[1]<<4)+(in_buffer[1]<<7))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<5)+(in_buffer[3]<<6))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<3)+(in_buffer[4]<<5))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<4)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<3)+(in_buffer[6]<<6))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<3))-(0+(in_buffer[8]<<4))-(0+(in_buffer[9]<<6)+(in_buffer[9]<<7))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<3)+(in_buffer[10]<<4))+(0+(in_buffer[11]<<4)+(in_buffer[11]<<5))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<1)+(in_buffer[12]<<4))-(0+(in_buffer[13]<<3)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<5))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<1)+(in_buffer[15]<<4))-(0+(in_buffer[16]<<3)+(in_buffer[16]<<4))+(0+(in_buffer[17]<<3))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<3)+(in_buffer[19]<<5))+(0-(in_buffer[20]<<0)-(in_buffer[20]<<2)+(in_buffer[20]<<4)+(in_buffer[20]<<5))+(0+(in_buffer[21]<<0)-(in_buffer[21]<<2)+(in_buffer[21]<<5))-(0+(in_buffer[22]<<1)+(in_buffer[22]<<3)+(in_buffer[22]<<4))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)+(in_buffer[23]<<5))-(0-(in_buffer[24]<<0)+(in_buffer[24]<<4)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<5))-(0-(in_buffer[1]<<0)+(in_buffer[1]<<3))-(0+(in_buffer[2]<<5))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<5))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<1))-(0-(in_buffer[6]<<1)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<3))+(0+(in_buffer[8]<<2))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2))-(0-(in_buffer[10]<<1)+(in_buffer[10]<<7))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<4))+(0+(in_buffer[12]<<3)+(in_buffer[12]<<5)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2)+(in_buffer[13]<<3))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<6))-(0+(in_buffer[15]<<0))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<2)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<1)+(in_buffer[17]<<3)+(in_buffer[17]<<6))+(0+(in_buffer[18]<<1)+(in_buffer[18]<<3)+(in_buffer[18]<<6))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<2)+(in_buffer[20]<<6))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<3))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)+(in_buffer[23]<<5))-(0-(in_buffer[24]<<0)-(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<4)+(in_buffer[0]<<7))-(0-(in_buffer[1]<<2)-(in_buffer[1]<<4)+(in_buffer[1]<<7))+(0+(in_buffer[2]<<3)+(in_buffer[2]<<5)+(in_buffer[2]<<6))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<6))-(0-(in_buffer[4]<<0)+(in_buffer[4]<<6))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<4))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<3)+(in_buffer[6]<<5))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<4))+(0-(in_buffer[8]<<2)+(in_buffer[8]<<6))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<5))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<5))-(0-(in_buffer[12]<<0)+(in_buffer[12]<<4))-(0+(in_buffer[13]<<0))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<1)+(in_buffer[14]<<5))+(0+(in_buffer[15]<<2)+(in_buffer[15]<<4))+(0+(in_buffer[16]<<1)+(in_buffer[16]<<3)+(in_buffer[16]<<6))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<3))-(0+(in_buffer[19]<<2)+(in_buffer[19]<<3))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<4)+(in_buffer[21]<<5))-(0+(in_buffer[22]<<2)+(in_buffer[22]<<3))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<3)+(in_buffer[23]<<5))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<4)+(in_buffer[0]<<7))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<3))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<1)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<3))-(0+(in_buffer[4]<<2)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<2)+(in_buffer[5]<<4)+(in_buffer[5]<<5))-(0+(in_buffer[7]<<4))-(0+(in_buffer[8]<<0)+(in_buffer[8]<<2))+(0-(in_buffer[9]<<0)+(in_buffer[9]<<4)+(in_buffer[9]<<5))-(0-(in_buffer[10]<<0)+(in_buffer[10]<<4)+(in_buffer[10]<<7))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<1)+(in_buffer[11]<<5))+(0-(in_buffer[12]<<1)+(in_buffer[12]<<7))-(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<6))-(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<5))+(0-(in_buffer[15]<<2)+(in_buffer[15]<<5)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<0)-(in_buffer[16]<<2)+(in_buffer[16]<<6))-(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<5))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<3)+(in_buffer[18]<<4))-(0-(in_buffer[19]<<0)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0-(in_buffer[21]<<1)-(in_buffer[21]<<3)+(in_buffer[21]<<6))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<3))-(0+(in_buffer[23]<<2)+(in_buffer[23]<<3))-(0-(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<4)+(in_buffer[24]<<7)+(in_buffer[24]<<8));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)-(in_buffer[0]<<4)+(in_buffer[0]<<6)+(in_buffer[0]<<7))+(0-(in_buffer[1]<<0)+(in_buffer[1]<<3)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<2)+(in_buffer[2]<<4))-(0-(in_buffer[3]<<2)+(in_buffer[3]<<5))+(0+(in_buffer[4]<<3)+(in_buffer[4]<<4))-(0-(in_buffer[5]<<2)-(in_buffer[5]<<4)+(in_buffer[5]<<8))+(0-(in_buffer[6]<<2)+(in_buffer[6]<<5))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<3))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<3)+(in_buffer[8]<<4))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<4)+(in_buffer[9]<<5))-(0+(in_buffer[10]<<4)+(in_buffer[10]<<6))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<3)+(in_buffer[11]<<6))-(0-(in_buffer[12]<<2)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<1)+(in_buffer[13]<<3)+(in_buffer[13]<<4))-(0-(in_buffer[14]<<0)+(in_buffer[14]<<3)+(in_buffer[14]<<4)+(in_buffer[14]<<7))+(0+(in_buffer[15]<<2)+(in_buffer[15]<<5))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<3))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<6))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<5)+(in_buffer[19]<<6))-(0-(in_buffer[20]<<2)+(in_buffer[20]<<4)+(in_buffer[20]<<5))+(0+(in_buffer[21]<<2)+(in_buffer[21]<<4))-(0-(in_buffer[22]<<2)+(in_buffer[22]<<4)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<0)-(in_buffer[23]<<3)+(in_buffer[23]<<6))-(0+(in_buffer[24]<<2)-(in_buffer[24]<<4)+(in_buffer[24]<<7));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight10;
assign in_buffer_weight10=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<5)+(in_buffer[0]<<6))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<4)+(in_buffer[1]<<5))-(0-(in_buffer[2]<<2)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<2)+(in_buffer[3]<<5))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<2)+(in_buffer[4]<<7))-(0+(in_buffer[5]<<4)+(in_buffer[5]<<5))-(0+(in_buffer[6]<<1)+(in_buffer[6]<<2))+(0+(in_buffer[7]<<4))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<1))+(0-(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<3))+(0+(in_buffer[10]<<4))+(0-(in_buffer[11]<<2)+(in_buffer[11]<<5)+(in_buffer[11]<<6))+(0+(in_buffer[12]<<0))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<4)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<3))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<5))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<2))-(0-(in_buffer[17]<<0)+(in_buffer[17]<<3)+(in_buffer[17]<<5))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<1)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<3)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<3)+(in_buffer[20]<<5))-(0+(in_buffer[21]<<1)+(in_buffer[21]<<3))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<6))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight11;
assign in_buffer_weight11=0-(0+(in_buffer[0]<<1)+(in_buffer[0]<<4)+(in_buffer[0]<<5))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<1))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<2)+(in_buffer[2]<<3))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<3))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<3))+(0+(in_buffer[5]<<1))+(0-(in_buffer[6]<<1)+(in_buffer[6]<<4))-(0-(in_buffer[7]<<1)-(in_buffer[7]<<3)+(in_buffer[7]<<5)+(in_buffer[7]<<6))+(0+(in_buffer[8]<<2)+(in_buffer[8]<<4)+(in_buffer[8]<<5))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<4))-(0+(in_buffer[10]<<4)+(in_buffer[10]<<5))-(0+(in_buffer[11]<<1)+(in_buffer[11]<<3))-(0-(in_buffer[12]<<3)+(in_buffer[12]<<5)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<1)+(in_buffer[13]<<2))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<4)+(in_buffer[14]<<5))+(0+(in_buffer[15]<<1)+(in_buffer[15]<<2)+(in_buffer[15]<<5)+(in_buffer[15]<<6))+(0+(in_buffer[16]<<4)+(in_buffer[16]<<5))+(0-(in_buffer[17]<<1)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<6))+(0-(in_buffer[19]<<3)+(in_buffer[19]<<6))-(0+(in_buffer[20]<<3)+(in_buffer[20]<<4))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<2)+(in_buffer[22]<<4))+(0-(in_buffer[23]<<2)+(in_buffer[23]<<5))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight12;
assign in_buffer_weight12=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<6))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<3)+(in_buffer[1]<<4)+(in_buffer[1]<<7))-(0+(in_buffer[2]<<3)+(in_buffer[2]<<6))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<4))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<3)+(in_buffer[4]<<4))+(0+(in_buffer[5]<<2)+(in_buffer[5]<<3))-(0-(in_buffer[6]<<1)+(in_buffer[6]<<4))+(0-(in_buffer[7]<<0)+(in_buffer[7]<<6))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<2)+(in_buffer[8]<<3))+(0-(in_buffer[9]<<1)+(in_buffer[9]<<5))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<6))-(0+(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<4)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<2)+(in_buffer[14]<<4))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<3))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<0)-(in_buffer[17]<<3)+(in_buffer[17]<<5)+(in_buffer[17]<<6))-(0+(in_buffer[18]<<2)+(in_buffer[18]<<3))-(0+(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<4)+(in_buffer[21]<<5))+(0-(in_buffer[22]<<2)+(in_buffer[22]<<6))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<5))+(0-(in_buffer[24]<<1)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight13;
assign in_buffer_weight13=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3))+(0+(in_buffer[1]<<0)-(in_buffer[1]<<2)+(in_buffer[1]<<6))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<3))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<2))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<2)+(in_buffer[4]<<6))-(0+(in_buffer[5]<<3))+(0+(in_buffer[6]<<0))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<4)+(in_buffer[7]<<6))-(0+(in_buffer[8]<<0))+(0-(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<3))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<2))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<4))+(0-(in_buffer[12]<<1)-(in_buffer[12]<<3)+(in_buffer[12]<<6))+(0+(in_buffer[13]<<3)+(in_buffer[13]<<4))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<4))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<3)+(in_buffer[15]<<4))+(0+(in_buffer[16]<<0))+(0-(in_buffer[17]<<2)+(in_buffer[17]<<6))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<4))+(0-(in_buffer[19]<<2)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<2))+(0+(in_buffer[21]<<2)+(in_buffer[21]<<4))-(0+(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<4)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<4))+(0+(in_buffer[24]<<0)-(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight14;
assign in_buffer_weight14=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<4))-(0+(in_buffer[1]<<1))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<3))-(0+(in_buffer[3]<<1))+(0+(in_buffer[4]<<1))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<1))+(0+(in_buffer[6]<<2)+(in_buffer[6]<<3))-(0+(in_buffer[7]<<1)+(in_buffer[7]<<4))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<1))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<1))+(0+(in_buffer[10]<<1)+(in_buffer[10]<<3))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<3))-(0+(in_buffer[12]<<3)+(in_buffer[12]<<4))+(0+(in_buffer[13]<<4))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<4))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<3)+(in_buffer[15]<<4))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<1)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<1)+(in_buffer[17]<<4))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<2))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<3))+(0+(in_buffer[21]<<1))-(0+(in_buffer[22]<<2)+(in_buffer[22]<<4))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<2))-(0-(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight15;
assign in_buffer_weight15=0-(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<3))+(0-(in_buffer[2]<<1)+(in_buffer[2]<<3)+(in_buffer[2]<<4))-(0-(in_buffer[3]<<1)+(in_buffer[3]<<3)+(in_buffer[3]<<4))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<3))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<3))+(0-(in_buffer[8]<<0)+(in_buffer[8]<<3)+(in_buffer[8]<<4))-(0-(in_buffer[9]<<1)+(in_buffer[9]<<4))-(0+(in_buffer[10]<<3)+(in_buffer[10]<<4))-(0-(in_buffer[11]<<0)+(in_buffer[11]<<3))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<2))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<1))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<4))-(0+(in_buffer[15]<<0))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<2))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<4))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<2))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<2))-(0+(in_buffer[22]<<3)+(in_buffer[22]<<4))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<2))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight16;
assign in_buffer_weight16=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<1)+(in_buffer[0]<<5)+(in_buffer[0]<<6))-(0+(in_buffer[1]<<0)-(in_buffer[1]<<3)+(in_buffer[1]<<5)+(in_buffer[1]<<6))-(0+(in_buffer[2]<<0)+(in_buffer[2]<<1)+(in_buffer[2]<<6))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<4)+(in_buffer[4]<<6))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<3))+(0+(in_buffer[6]<<2)+(in_buffer[6]<<4))-(0+(in_buffer[7]<<1)+(in_buffer[7]<<3))+(0+(in_buffer[8]<<5))+(0+(in_buffer[9]<<2)+(in_buffer[9]<<6))+(0-(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<4)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<5)+(in_buffer[11]<<6))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<3))+(0+(in_buffer[13]<<2)+(in_buffer[13]<<3))-(0+(in_buffer[14]<<3))-(0+(in_buffer[15]<<6))-(0+(in_buffer[16]<<0)-(in_buffer[16]<<3)+(in_buffer[16]<<6))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<5))+(0+(in_buffer[18]<<1)+(in_buffer[18]<<2))-(0+(in_buffer[19]<<0)+(in_buffer[19]<<1)+(in_buffer[19]<<4))+(0-(in_buffer[20]<<1)+(in_buffer[20]<<4)+(in_buffer[20]<<5))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<3))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<3))+(0+(in_buffer[24]<<3)+(in_buffer[24]<<4));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight17;
assign in_buffer_weight17=0-(0+(in_buffer[0]<<2)-(in_buffer[0]<<4)+(in_buffer[0]<<7))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<3)+(in_buffer[2]<<4))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<1))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<1))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<4)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<5))+(0-(in_buffer[7]<<0)+(in_buffer[7]<<5))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<5))-(0+(in_buffer[9]<<0))+(0-(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<6))+(0+(in_buffer[12]<<1)+(in_buffer[12]<<4))-(0+(in_buffer[13]<<1)+(in_buffer[13]<<3))-(0-(in_buffer[14]<<3)+(in_buffer[14]<<6))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<4)+(in_buffer[15]<<5))-(0-(in_buffer[16]<<1)+(in_buffer[16]<<4))+(0-(in_buffer[17]<<1)+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<5))-(0+(in_buffer[19]<<1)+(in_buffer[19]<<4)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<6))-(0+(in_buffer[21]<<1)+(in_buffer[21]<<3))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<2)+(in_buffer[22]<<6))+(0+(in_buffer[23]<<3)+(in_buffer[23]<<7))+(0-(in_buffer[24]<<1)+(in_buffer[24]<<5)+(in_buffer[24]<<7));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight18;
assign in_buffer_weight18=0-(0-(in_buffer[0]<<0)-(in_buffer[0]<<3)+(in_buffer[0]<<6))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<1)+(in_buffer[1]<<4)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<0)-(in_buffer[2]<<3)+(in_buffer[2]<<5)+(in_buffer[2]<<6))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<4))-(0+(in_buffer[4]<<1)-(in_buffer[4]<<4)+(in_buffer[4]<<8))+(0+(in_buffer[5]<<2)+(in_buffer[5]<<4)+(in_buffer[5]<<5))+(0+(in_buffer[6]<<2)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<5))+(0-(in_buffer[8]<<2)+(in_buffer[8]<<5))-(0+(in_buffer[9]<<4))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<1)+(in_buffer[11]<<4)+(in_buffer[11]<<5))-(0-(in_buffer[12]<<2)+(in_buffer[12]<<6))+(0-(in_buffer[13]<<1)+(in_buffer[13]<<4)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<5))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3))-(0-(in_buffer[16]<<1)+(in_buffer[16]<<4))+(0+(in_buffer[17]<<2)+(in_buffer[17]<<4))-(0-(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<3))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<2))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<1)+(in_buffer[20]<<5))+(0-(in_buffer[21]<<0)-(in_buffer[21]<<2)+(in_buffer[21]<<5))+(0-(in_buffer[22]<<0)+(in_buffer[22]<<6))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)+(in_buffer[23]<<4))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight19;
assign in_buffer_weight19=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<1)+(in_buffer[0]<<7))+(0-(in_buffer[1]<<1)+(in_buffer[1]<<4)+(in_buffer[1]<<5))-(0-(in_buffer[2]<<1)+(in_buffer[2]<<4))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<3))+(0-(in_buffer[4]<<1)+(in_buffer[4]<<5))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3))-(0-(in_buffer[6]<<0)-(in_buffer[6]<<2)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<1)+(in_buffer[7]<<3)+(in_buffer[7]<<4))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<3)+(in_buffer[8]<<4))-(0-(in_buffer[9]<<0)+(in_buffer[9]<<3)+(in_buffer[9]<<4))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<5))+(0+(in_buffer[12]<<1)+(in_buffer[12]<<5))+(0+(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<4)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<5))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<1)+(in_buffer[15]<<6))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<4)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<2))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<5)+(in_buffer[19]<<6))+(0+(in_buffer[20]<<0))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<5))-(0-(in_buffer[22]<<2)+(in_buffer[22]<<4)+(in_buffer[22]<<5))-(0-(in_buffer[23]<<2)+(in_buffer[23]<<6)+(in_buffer[23]<<8))-(0-(in_buffer[24]<<0)-(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight20;
assign in_buffer_weight20=0-(0+(in_buffer[0]<<4))+(0+(in_buffer[1]<<2)+(in_buffer[1]<<4)+(in_buffer[1]<<5))+(0-(in_buffer[2]<<0)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<6))-(0-(in_buffer[4]<<0)+(in_buffer[4]<<4)+(in_buffer[4]<<5))+(0+(in_buffer[5]<<0)+(in_buffer[5]<<1))-(0+(in_buffer[6]<<5))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<4))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<1)+(in_buffer[8]<<4))-(0-(in_buffer[9]<<0)+(in_buffer[9]<<3))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<3))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<6))+(0+(in_buffer[13]<<0)+(in_buffer[13]<<6))+(0+(in_buffer[14]<<5))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<2))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<3)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<6))+(0-(in_buffer[18]<<0)+(in_buffer[18]<<4)+(in_buffer[18]<<5))-(0-(in_buffer[19]<<0)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<3))+(0+(in_buffer[21]<<3))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<2)+(in_buffer[22]<<4))+(0+(in_buffer[23]<<3)+(in_buffer[23]<<4))-(0-(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<5)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight21;
assign in_buffer_weight21=0-(0+(in_buffer[0]<<1)+(in_buffer[0]<<4)-(in_buffer[0]<<6)+(in_buffer[0]<<9))-(0+(in_buffer[1]<<2)+(in_buffer[1]<<5))+(0-(in_buffer[2]<<3)+(in_buffer[2]<<5)+(in_buffer[2]<<6))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<1)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<1)+(in_buffer[5]<<3)+(in_buffer[5]<<4)+(in_buffer[5]<<7))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<4)+(in_buffer[6]<<5))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<5))+(0+(in_buffer[8]<<2)+(in_buffer[8]<<4))+(0+(in_buffer[9]<<2)+(in_buffer[9]<<6))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<1))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<6))+(0-(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<3))+(0+(in_buffer[13]<<1))+(0-(in_buffer[14]<<1)+(in_buffer[14]<<5))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<5)+(in_buffer[15]<<6))-(0+(in_buffer[17]<<1)+(in_buffer[17]<<4))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<3))-(0+(in_buffer[19]<<2)+(in_buffer[19]<<5)+(in_buffer[19]<<6))-(0-(in_buffer[21]<<1)+(in_buffer[21]<<4))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<2))-(0-(in_buffer[23]<<0)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<1)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight22;
assign in_buffer_weight22=0-(0-(in_buffer[0]<<1)+(in_buffer[0]<<5)+(in_buffer[0]<<6))-(0-(in_buffer[1]<<1)+(in_buffer[1]<<4))-(0-(in_buffer[2]<<0)+(in_buffer[2]<<3)+(in_buffer[2]<<4))+(0+(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<5))-(0+(in_buffer[4]<<3))+(0+(in_buffer[5]<<4)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<2)+(in_buffer[6]<<3))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<4))+(0+(in_buffer[8]<<1))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<3)+(in_buffer[9]<<4))-(0-(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<5)+(in_buffer[10]<<6))-(0-(in_buffer[11]<<1)-(in_buffer[11]<<3)+(in_buffer[11]<<5)+(in_buffer[11]<<6))+(0-(in_buffer[12]<<1)+(in_buffer[12]<<5)+(in_buffer[12]<<6))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<4))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<3))-(0+(in_buffer[15]<<2)+(in_buffer[15]<<4))+(0+(in_buffer[16]<<1)+(in_buffer[16]<<4)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<3))-(0+(in_buffer[18]<<3))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<2)+(in_buffer[19]<<4))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<4))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<3))-(0+(in_buffer[22]<<1)+(in_buffer[22]<<4))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<2))+(0-(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight23;
assign in_buffer_weight23=0-(0+(in_buffer[0]<<4))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<1)+(in_buffer[1]<<5))-(0-(in_buffer[2]<<0)+(in_buffer[2]<<3)+(in_buffer[2]<<4))+(0+(in_buffer[3]<<2))+(0+(in_buffer[4]<<0)-(in_buffer[4]<<3)+(in_buffer[4]<<5)+(in_buffer[4]<<6))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3))-(0-(in_buffer[6]<<0)+(in_buffer[6]<<3))+(0+(in_buffer[7]<<2)+(in_buffer[7]<<3))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<5))-(0-(in_buffer[9]<<0)+(in_buffer[9]<<4)+(in_buffer[9]<<5))-(0+(in_buffer[10]<<0))-(0+(in_buffer[11]<<1)+(in_buffer[11]<<2)+(in_buffer[11]<<5))-(0+(in_buffer[12]<<1)+(in_buffer[12]<<3)+(in_buffer[12]<<4))+(0+(in_buffer[13]<<1)-(in_buffer[13]<<3)+(in_buffer[13]<<6))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<4)+(in_buffer[14]<<5))+(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<7))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<6))-(0+(in_buffer[17]<<3)+(in_buffer[17]<<5))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<1)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<3))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<3)+(in_buffer[20]<<7))-(0+(in_buffer[21]<<6))+(0+(in_buffer[22]<<2)+(in_buffer[22]<<4)+(in_buffer[22]<<5))+(0-(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<4)+(in_buffer[23]<<5))-(0-(in_buffer[24]<<2)+(in_buffer[24]<<5)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight24;
assign in_buffer_weight24=0+(0+(in_buffer[0]<<2)+(in_buffer[0]<<4)+(in_buffer[0]<<5))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<2))-(0-(in_buffer[2]<<0)+(in_buffer[2]<<4))-(0-(in_buffer[3]<<0)+(in_buffer[3]<<3))-(0+(in_buffer[4]<<1)+(in_buffer[4]<<4))+(0-(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<4)+(in_buffer[5]<<5))+(0+(in_buffer[6]<<1)+(in_buffer[6]<<3))-(0+(in_buffer[7]<<4)+(in_buffer[7]<<5))+(0-(in_buffer[8]<<1)+(in_buffer[8]<<5))+(0-(in_buffer[9]<<1)+(in_buffer[9]<<5))+(0+(in_buffer[10]<<3)+(in_buffer[10]<<4))-(0+(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<4))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<1)+(in_buffer[12]<<5))+(0+(in_buffer[13]<<0))+(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<6))-(0-(in_buffer[15]<<1)-(in_buffer[15]<<3)+(in_buffer[15]<<6))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<4)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<1))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<1)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<4))-(0+(in_buffer[20]<<4)+(in_buffer[20]<<6))-(0+(in_buffer[21]<<1)+(in_buffer[21]<<4))+(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)+(in_buffer[23]<<4))-(0-(in_buffer[24]<<1)-(in_buffer[24]<<3)+(in_buffer[24]<<7));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight25;
assign in_buffer_weight25=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<1)+(in_buffer[0]<<6)+(in_buffer[0]<<7))+(0+(in_buffer[1]<<0)-(in_buffer[1]<<2)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<1)-(in_buffer[2]<<3)+(in_buffer[2]<<5)+(in_buffer[2]<<6))-(0+(in_buffer[3]<<4)+(in_buffer[3]<<6))+(0+(in_buffer[4]<<4))-(0-(in_buffer[5]<<2)+(in_buffer[5]<<5)+(in_buffer[5]<<7))-(0-(in_buffer[6]<<0)-(in_buffer[6]<<3)+(in_buffer[6]<<7))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<4))+(0-(in_buffer[8]<<1)+(in_buffer[8]<<4))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<1)+(in_buffer[9]<<6))-(0+(in_buffer[10]<<2)+(in_buffer[10]<<4))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<4)+(in_buffer[11]<<5))-(0-(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<5))-(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<5))-(0-(in_buffer[14]<<1)+(in_buffer[14]<<6))+(0+(in_buffer[15]<<0)-(in_buffer[15]<<3)+(in_buffer[15]<<5)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<3)+(in_buffer[16]<<5))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<6))+(0+(in_buffer[19]<<0)-(in_buffer[19]<<2)+(in_buffer[19]<<4)+(in_buffer[19]<<5))-(0-(in_buffer[20]<<1)+(in_buffer[20]<<5))-(0+(in_buffer[21]<<0))+(0+(in_buffer[22]<<3)+(in_buffer[22]<<4))-(0-(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<4))+(0+(in_buffer[24]<<1)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight26;
assign in_buffer_weight26=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<5))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<1)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<2))-(0+(in_buffer[3]<<0))-(0-(in_buffer[4]<<0)+(in_buffer[4]<<3)+(in_buffer[4]<<5))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<4)+(in_buffer[6]<<5))+(0-(in_buffer[7]<<2)+(in_buffer[7]<<6))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<3))+(0+(in_buffer[9]<<0))-(0-(in_buffer[10]<<0)+(in_buffer[10]<<3)+(in_buffer[10]<<5))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<7))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<1)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2)+(in_buffer[13]<<3))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<4))+(0+(in_buffer[15]<<2)+(in_buffer[15]<<6))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<4)+(in_buffer[17]<<6))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<3)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<2)+(in_buffer[19]<<6))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<2)+(in_buffer[20]<<4)+(in_buffer[20]<<5))-(0+(in_buffer[21]<<4))+(0+(in_buffer[22]<<5))-(0+(in_buffer[23]<<5))-(0-(in_buffer[24]<<3)-(in_buffer[24]<<5)+(in_buffer[24]<<7)+(in_buffer[24]<<8));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight27;
assign in_buffer_weight27=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3))+(0-(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<3))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<2)+(in_buffer[2]<<3)+(in_buffer[2]<<6))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<3)+(in_buffer[3]<<4))-(0-(in_buffer[4]<<0)-(in_buffer[4]<<2)+(in_buffer[4]<<4)+(in_buffer[4]<<5))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<4))+(0-(in_buffer[6]<<1)+(in_buffer[6]<<3)+(in_buffer[6]<<4))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<4))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<4)+(in_buffer[8]<<5))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<4))+(0+(in_buffer[10]<<1)+(in_buffer[10]<<2))+(0+(in_buffer[11]<<0)-(in_buffer[11]<<3)+(in_buffer[11]<<6))-(0-(in_buffer[12]<<1)+(in_buffer[12]<<4))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<3)+(in_buffer[13]<<4))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<2))-(0+(in_buffer[15]<<1)+(in_buffer[15]<<3)+(in_buffer[15]<<5))+(0-(in_buffer[16]<<1)+(in_buffer[16]<<6))+(0+(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<4))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<4))+(0-(in_buffer[21]<<1)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<5))-(0-(in_buffer[23]<<0)-(in_buffer[23]<<3)+(in_buffer[23]<<5)+(in_buffer[23]<<6))-(0-(in_buffer[24]<<2)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight28;
assign in_buffer_weight28=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<4))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<2)+(in_buffer[1]<<5))-(0+(in_buffer[2]<<1))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<2)+(in_buffer[3]<<5))+(0-(in_buffer[4]<<1)+(in_buffer[4]<<3)+(in_buffer[4]<<4))+(0-(in_buffer[5]<<1)+(in_buffer[5]<<4)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<2)+(in_buffer[6]<<4))+(0+(in_buffer[7]<<3))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<3))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<3)+(in_buffer[9]<<4))-(0-(in_buffer[10]<<2)-(in_buffer[10]<<4)+(in_buffer[10]<<7))-(0-(in_buffer[11]<<1)+(in_buffer[11]<<6))+(0-(in_buffer[12]<<0)+(in_buffer[12]<<3))+(0+(in_buffer[13]<<1)+(in_buffer[13]<<4)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<5))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<1)-(in_buffer[15]<<4)+(in_buffer[15]<<7)+(in_buffer[15]<<8))+(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<3))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<6))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<1)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)-(in_buffer[20]<<5)+(in_buffer[20]<<7)+(in_buffer[20]<<8))-(0-(in_buffer[21]<<3)+(in_buffer[21]<<6))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<6))+(0+(in_buffer[23]<<0))-(0+(in_buffer[24]<<1)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight29;
assign in_buffer_weight29=0-(0-(in_buffer[0]<<2)+(in_buffer[0]<<5))-(0-(in_buffer[1]<<1)+(in_buffer[1]<<4))-(0-(in_buffer[2]<<1)+(in_buffer[2]<<4)+(in_buffer[2]<<5))+(0-(in_buffer[3]<<1)+(in_buffer[3]<<5)+(in_buffer[3]<<6))-(0-(in_buffer[4]<<0)+(in_buffer[4]<<3)+(in_buffer[4]<<4))-(0+(in_buffer[5]<<1))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<2))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<2)+(in_buffer[7]<<4))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<5))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<4))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<2))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<4)+(in_buffer[11]<<5))-(0-(in_buffer[12]<<0)+(in_buffer[12]<<3))+(0+(in_buffer[13]<<0)+(in_buffer[13]<<1)+(in_buffer[13]<<4)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<6))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<5)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<3)+(in_buffer[16]<<6))+(0-(in_buffer[17]<<1)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<1)+(in_buffer[18]<<3))-(0-(in_buffer[19]<<0)-(in_buffer[19]<<3)+(in_buffer[19]<<5)+(in_buffer[19]<<6))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<2)+(in_buffer[20]<<5)+(in_buffer[20]<<6))-(0-(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<8))+(0-(in_buffer[22]<<0)+(in_buffer[22]<<2)+(in_buffer[22]<<3)+(in_buffer[22]<<6))+(0-(in_buffer[23]<<1)+(in_buffer[23]<<5))+(0+(in_buffer[24]<<1)+(in_buffer[24]<<2)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight30;
assign in_buffer_weight30=0+(0+(in_buffer[0]<<1)+(in_buffer[0]<<3)+(in_buffer[0]<<4))-(0+(in_buffer[1]<<3))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<3)+(in_buffer[2]<<4))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<1)-(in_buffer[3]<<4)+(in_buffer[3]<<7))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<4)+(in_buffer[4]<<7))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<4))+(0+(in_buffer[6]<<1))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<4))-(0+(in_buffer[8]<<0)+(in_buffer[8]<<7))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<3)+(in_buffer[9]<<6)+(in_buffer[9]<<7))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<2))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3))-(0-(in_buffer[12]<<0)+(in_buffer[12]<<4))+(0-(in_buffer[13]<<0)+(in_buffer[13]<<3)+(in_buffer[13]<<6))+(0-(in_buffer[14]<<1)+(in_buffer[14]<<4))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<4))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<3))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<3)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<5))+(0-(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<4))+(0-(in_buffer[20]<<1)+(in_buffer[20]<<4))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<3)+(in_buffer[21]<<4))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<3)+(in_buffer[22]<<5))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<4)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight31;
assign in_buffer_weight31=0-(0+(in_buffer[0]<<4))-(0-(in_buffer[1]<<2)+(in_buffer[1]<<5))-(0-(in_buffer[2]<<2)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<2)+(in_buffer[3]<<4))-(0+(in_buffer[4]<<1)+(in_buffer[4]<<2))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<4))-(0+(in_buffer[6]<<1)+(in_buffer[6]<<2))+(0+(in_buffer[7]<<0))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<3)+(in_buffer[8]<<4))+(0+(in_buffer[9]<<1))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<2))-(0+(in_buffer[11]<<1)+(in_buffer[11]<<2))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<4))-(0+(in_buffer[14]<<1)+(in_buffer[14]<<3)+(in_buffer[14]<<4))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<3)+(in_buffer[17]<<4))+(0-(in_buffer[18]<<0)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<2)+(in_buffer[19]<<4))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<2))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<4))-(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<4))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<4));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight32;
assign in_buffer_weight32=0-(0-(in_buffer[0]<<0)-(in_buffer[0]<<3)+(in_buffer[0]<<7)+(in_buffer[0]<<8))-(0+(in_buffer[1]<<4)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<2)+(in_buffer[2]<<6))+(0-(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<5))-(0+(in_buffer[4]<<2)+(in_buffer[4]<<3))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<1)+(in_buffer[6]<<4)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<1))-(0+(in_buffer[8]<<4)+(in_buffer[8]<<5))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<4)+(in_buffer[9]<<5))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<3)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<2))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<3)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<1)-(in_buffer[13]<<3)+(in_buffer[13]<<5)+(in_buffer[13]<<6))-(0-(in_buffer[14]<<4)+(in_buffer[14]<<7))-(0+(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<4)+(in_buffer[15]<<5))+(0+(in_buffer[16]<<2))-(0+(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<3))+(0-(in_buffer[19]<<0)-(in_buffer[19]<<2)-(in_buffer[19]<<4)+(in_buffer[19]<<7))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<2)+(in_buffer[20]<<6))-(0-(in_buffer[21]<<2)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<3)+(in_buffer[22]<<5))+(0-(in_buffer[23]<<1)-(in_buffer[23]<<3)+(in_buffer[23]<<6))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight33;
assign in_buffer_weight33=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<1)-(in_buffer[0]<<4)+(in_buffer[0]<<6)+(in_buffer[0]<<7))-(0+(in_buffer[1]<<1)-(in_buffer[1]<<3)+(in_buffer[1]<<7))-(0+(in_buffer[2]<<0)+(in_buffer[2]<<1)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<4))+(0-(in_buffer[4]<<1)+(in_buffer[4]<<4)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<1)-(in_buffer[5]<<3)-(in_buffer[5]<<5)+(in_buffer[5]<<7)+(in_buffer[5]<<8))-(0+(in_buffer[6]<<5)+(in_buffer[6]<<6))+(0-(in_buffer[7]<<1)-(in_buffer[7]<<3)+(in_buffer[7]<<5)+(in_buffer[7]<<6))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<6))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<3)+(in_buffer[9]<<4))-(0+(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<6))-(0+(in_buffer[11]<<3))+(0-(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<5)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<3)+(in_buffer[13]<<4))-(0+(in_buffer[14]<<0)-(in_buffer[14]<<3)+(in_buffer[14]<<5)+(in_buffer[14]<<6))-(0-(in_buffer[15]<<1)+(in_buffer[15]<<3)+(in_buffer[15]<<4))-(0-(in_buffer[16]<<2)+(in_buffer[16]<<5))+(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0-(in_buffer[18]<<0)+(in_buffer[18]<<3)+(in_buffer[18]<<4))+(0-(in_buffer[19]<<1)+(in_buffer[19]<<4)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)-(in_buffer[20]<<4)+(in_buffer[20]<<7))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<3))+(0+(in_buffer[22]<<0))+(0-(in_buffer[23]<<1)+(in_buffer[23]<<4))+(0+(in_buffer[24]<<0));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight34;
assign in_buffer_weight34=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<5)+(in_buffer[1]<<6))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<3))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<2)+(in_buffer[3]<<5))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<3)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<1)-(in_buffer[5]<<3)+(in_buffer[5]<<5)+(in_buffer[5]<<6))+(0+(in_buffer[6]<<0))-(0+(in_buffer[7]<<5))-(0+(in_buffer[8]<<1))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<5))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<3))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<4)+(in_buffer[11]<<5))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<2))+(0+(in_buffer[13]<<2)+(in_buffer[13]<<4))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<5))-(0-(in_buffer[15]<<1)+(in_buffer[15]<<7))+(0+(in_buffer[16]<<1)+(in_buffer[16]<<2)+(in_buffer[16]<<6))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<4)+(in_buffer[17]<<5))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<4))-(0+(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<2))-(0+(in_buffer[21]<<1)+(in_buffer[21]<<5)+(in_buffer[21]<<6))-(0-(in_buffer[22]<<0)+(in_buffer[22]<<4)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<1)-(in_buffer[23]<<3)+(in_buffer[23]<<6))+(0-(in_buffer[24]<<1)-(in_buffer[24]<<3)+(in_buffer[24]<<6)+(in_buffer[24]<<7));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight35;
assign in_buffer_weight35=0+(0+(in_buffer[0]<<2)+(in_buffer[0]<<6))+(0+(in_buffer[1]<<1))-(0+(in_buffer[2]<<0))-(0-(in_buffer[3]<<0)+(in_buffer[3]<<4)+(in_buffer[3]<<5))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<2))-(0+(in_buffer[5]<<2)+(in_buffer[5]<<5))+(0-(in_buffer[6]<<1)+(in_buffer[6]<<5))+(0+(in_buffer[7]<<2))+(0-(in_buffer[8]<<2)+(in_buffer[8]<<4)+(in_buffer[8]<<5))+(0+(in_buffer[9]<<0)-(in_buffer[9]<<3)+(in_buffer[9]<<5)+(in_buffer[9]<<6))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<3))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<4))+(0+(in_buffer[12]<<2)+(in_buffer[12]<<3))-(0-(in_buffer[13]<<1)+(in_buffer[13]<<3)+(in_buffer[13]<<4))-(0-(in_buffer[14]<<1)+(in_buffer[14]<<4)+(in_buffer[14]<<5))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<3)+(in_buffer[16]<<4))+(0+(in_buffer[17]<<5))-(0-(in_buffer[18]<<0)+(in_buffer[18]<<6))+(0+(in_buffer[19]<<0)-(in_buffer[19]<<2)+(in_buffer[19]<<4)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0-(in_buffer[21]<<2)+(in_buffer[21]<<6))-(0+(in_buffer[23]<<1)+(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<7)+(in_buffer[23]<<8))+(0+(in_buffer[24]<<0)-(in_buffer[24]<<4)+(in_buffer[24]<<7));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight36;
assign in_buffer_weight36=0-(0+(in_buffer[0]<<5))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<3))+(0+(in_buffer[2]<<4))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<2))+(0+(in_buffer[4]<<2)+(in_buffer[4]<<5))+(0-(in_buffer[5]<<1)+(in_buffer[5]<<5)+(in_buffer[5]<<7))+(0-(in_buffer[6]<<2)+(in_buffer[6]<<5)+(in_buffer[6]<<6))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<5))+(0+(in_buffer[8]<<0))-(0-(in_buffer[9]<<1)+(in_buffer[9]<<5))-(0-(in_buffer[10]<<3)+(in_buffer[10]<<6)+(in_buffer[10]<<7))-(0+(in_buffer[11]<<0)-(in_buffer[11]<<4)+(in_buffer[11]<<7))+(0+(in_buffer[12]<<6))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<1)+(in_buffer[14]<<5))+(0-(in_buffer[15]<<3)+(in_buffer[15]<<6))+(0-(in_buffer[16]<<1)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<1)+(in_buffer[18]<<3))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<5))+(0-(in_buffer[20]<<0)+(in_buffer[20]<<4)+(in_buffer[20]<<6))+(0+(in_buffer[21]<<2)+(in_buffer[21]<<3)+(in_buffer[21]<<6))+(0-(in_buffer[22]<<0)+(in_buffer[22]<<3))-(0+(in_buffer[23]<<1)+(in_buffer[23]<<3))+(0+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight37;
assign in_buffer_weight37=0+(0+(in_buffer[0]<<5)+(in_buffer[0]<<6))+(0-(in_buffer[1]<<1)+(in_buffer[1]<<5))-(0-(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<5))-(0-(in_buffer[3]<<0)+(in_buffer[3]<<4))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<5))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<2))+(0+(in_buffer[6]<<2)+(in_buffer[6]<<3)+(in_buffer[6]<<6))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<7))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<5))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<1)+(in_buffer[9]<<5))+(0-(in_buffer[10]<<1)+(in_buffer[10]<<4))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<4)+(in_buffer[11]<<6))+(0-(in_buffer[12]<<0)+(in_buffer[12]<<3)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<1)+(in_buffer[13]<<2))+(0+(in_buffer[14]<<1)+(in_buffer[14]<<3)+(in_buffer[14]<<4))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<3)+(in_buffer[15]<<5))-(0+(in_buffer[16]<<3)+(in_buffer[16]<<5))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0-(in_buffer[18]<<1)+(in_buffer[18]<<4))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<2)+(in_buffer[19]<<3))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<3)+(in_buffer[20]<<5)+(in_buffer[20]<<6))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<4))+(0-(in_buffer[22]<<1)+(in_buffer[22]<<3)+(in_buffer[22]<<4))-(0+(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<4))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight38;
assign in_buffer_weight38=0+(0-(in_buffer[0]<<3)+(in_buffer[0]<<5)+(in_buffer[0]<<6))+(0+(in_buffer[1]<<0)-(in_buffer[1]<<2)+(in_buffer[1]<<4)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<1)+(in_buffer[2]<<4)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<3))+(0-(in_buffer[4]<<0)+(in_buffer[4]<<4))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<1)+(in_buffer[5]<<4)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<4)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<4)+(in_buffer[7]<<6))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<5))-(0-(in_buffer[9]<<1)-(in_buffer[9]<<3)+(in_buffer[9]<<6))+(0-(in_buffer[10]<<0)+(in_buffer[10]<<3))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<6))+(0+(in_buffer[12]<<1)+(in_buffer[12]<<3)+(in_buffer[12]<<6))+(0+(in_buffer[13]<<3)+(in_buffer[13]<<4))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2))+(0+(in_buffer[15]<<2))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<3))-(0+(in_buffer[17]<<3)+(in_buffer[17]<<6))+(0+(in_buffer[18]<<2)+(in_buffer[18]<<5))+(0-(in_buffer[19]<<2)+(in_buffer[19]<<6))-(0-(in_buffer[20]<<3)+(in_buffer[20]<<5)+(in_buffer[20]<<6))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<5))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<1)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<1)+(in_buffer[23]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight39;
assign in_buffer_weight39=0+(0+(in_buffer[0]<<3))+(0-(in_buffer[1]<<2)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<2))+(0+(in_buffer[3]<<2)+(in_buffer[3]<<4))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<3)+(in_buffer[4]<<5))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<3))-(0+(in_buffer[6]<<0)-(in_buffer[6]<<2)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<1))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<4))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<2)+(in_buffer[9]<<5))-(0-(in_buffer[10]<<2)+(in_buffer[10]<<4)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<6))+(0-(in_buffer[12]<<0)-(in_buffer[12]<<3)+(in_buffer[12]<<6))-(0+(in_buffer[14]<<0))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<1)+(in_buffer[16]<<5)+(in_buffer[16]<<7))-(0-(in_buffer[17]<<0)+(in_buffer[17]<<5))+(0+(in_buffer[18]<<2)+(in_buffer[18]<<3))+(0-(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<4))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<4)+(in_buffer[20]<<6))+(0+(in_buffer[21]<<5)+(in_buffer[21]<<6))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<3))-(0-(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<4))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight40;
assign in_buffer_weight40=0-(0+(in_buffer[0]<<2)+(in_buffer[0]<<3))+(0-(in_buffer[1]<<0)+(in_buffer[1]<<3))+(0-(in_buffer[2]<<0)+(in_buffer[2]<<3))+(0-(in_buffer[3]<<0)+(in_buffer[3]<<3))+(0+(in_buffer[5]<<0)+(in_buffer[5]<<3))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<2))+(0+(in_buffer[7]<<1))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<2))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<3)+(in_buffer[9]<<4))-(0-(in_buffer[10]<<1)+(in_buffer[10]<<3)+(in_buffer[10]<<4))-(0-(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<4))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<2))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<2)+(in_buffer[13]<<3))+(0-(in_buffer[14]<<1)+(in_buffer[14]<<4))+(0+(in_buffer[16]<<0)+(in_buffer[16]<<1))-(0-(in_buffer[17]<<1)+(in_buffer[17]<<3)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<3))-(0+(in_buffer[19]<<0)+(in_buffer[19]<<3)+(in_buffer[19]<<4))-(0-(in_buffer[20]<<0)+(in_buffer[20]<<3)+(in_buffer[20]<<4))-(0+(in_buffer[21]<<2)+(in_buffer[21]<<4))-(0+(in_buffer[22]<<4))-(0+(in_buffer[23]<<4))-(0+(in_buffer[24]<<1)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight41;
assign in_buffer_weight41=0+(0-(in_buffer[0]<<3)+(in_buffer[0]<<6))+(0-(in_buffer[1]<<0)-(in_buffer[1]<<2)+(in_buffer[1]<<5))-(0+(in_buffer[2]<<4)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<4))+(0+(in_buffer[4]<<0)-(in_buffer[4]<<3)+(in_buffer[4]<<5)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<4))+(0-(in_buffer[6]<<2)+(in_buffer[6]<<5))+(0-(in_buffer[7]<<0)+(in_buffer[7]<<2)+(in_buffer[7]<<3))+(0+(in_buffer[8]<<3)+(in_buffer[8]<<4))-(0+(in_buffer[9]<<2)+(in_buffer[9]<<6))+(0-(in_buffer[10]<<2)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<6))-(0-(in_buffer[12]<<2)+(in_buffer[12]<<6))+(0+(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<5)+(in_buffer[13]<<6))+(0+(in_buffer[14]<<2))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<1)+(in_buffer[15]<<4))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<3)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<4))+(0+(in_buffer[18]<<5))-(0-(in_buffer[19]<<1)+(in_buffer[19]<<4)+(in_buffer[19]<<6))-(0-(in_buffer[20]<<3)+(in_buffer[20]<<5)+(in_buffer[20]<<6))-(0+(in_buffer[21]<<2)+(in_buffer[21]<<3)+(in_buffer[21]<<6))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<3)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<4));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight42;
assign in_buffer_weight42=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<5))+(0-(in_buffer[1]<<1)+(in_buffer[1]<<5))-(0+(in_buffer[2]<<2))+(0-(in_buffer[3]<<0)+(in_buffer[3]<<4)+(in_buffer[3]<<6))-(0+(in_buffer[4]<<1)+(in_buffer[4]<<2)+(in_buffer[4]<<5))-(0-(in_buffer[5]<<0)-(in_buffer[5]<<3)+(in_buffer[5]<<6))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<1)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<1)+(in_buffer[7]<<4)+(in_buffer[7]<<5))+(0-(in_buffer[8]<<0)+(in_buffer[8]<<7))+(0+(in_buffer[9]<<2)+(in_buffer[9]<<3))+(0-(in_buffer[10]<<1)+(in_buffer[10]<<4))-(0+(in_buffer[11]<<2))-(0+(in_buffer[12]<<4)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<4))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<6))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<3)+(in_buffer[15]<<4))-(0+(in_buffer[16]<<0)-(in_buffer[16]<<2)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<3))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<3)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<2)+(in_buffer[19]<<4))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0+(in_buffer[21]<<5))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<3)+(in_buffer[22]<<4))-(0+(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<6))+(0-(in_buffer[24]<<2)+(in_buffer[24]<<4)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight43;
assign in_buffer_weight43=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<4)+(in_buffer[0]<<6))+(0+(in_buffer[1]<<0)-(in_buffer[1]<<2)-(in_buffer[1]<<4)+(in_buffer[1]<<7))+(0+(in_buffer[2]<<0))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<1)+(in_buffer[3]<<4))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<5)+(in_buffer[4]<<6))+(0+(in_buffer[5]<<1)+(in_buffer[5]<<4)+(in_buffer[5]<<6))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<3)+(in_buffer[6]<<4))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<2)+(in_buffer[7]<<4))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<6))-(0-(in_buffer[9]<<2)+(in_buffer[9]<<7))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<4))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<3))-(0+(in_buffer[12]<<1)+(in_buffer[12]<<2)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<0))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<3)+(in_buffer[14]<<5))-(0-(in_buffer[15]<<1)+(in_buffer[15]<<7))-(0-(in_buffer[16]<<1)+(in_buffer[16]<<4)+(in_buffer[16]<<6))+(0+(in_buffer[17]<<1))+(0+(in_buffer[18]<<1)+(in_buffer[18]<<3)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<5))+(0-(in_buffer[20]<<0)-(in_buffer[20]<<3)+(in_buffer[20]<<8))+(0+(in_buffer[21]<<2)+(in_buffer[21]<<4)+(in_buffer[21]<<6))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<1)+(in_buffer[22]<<5))+(0+(in_buffer[23]<<2)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight44;
assign in_buffer_weight44=0+(0+(in_buffer[0]<<0)-(in_buffer[0]<<2)+(in_buffer[0]<<5))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<3)+(in_buffer[1]<<6))+(0+(in_buffer[2]<<2)+(in_buffer[2]<<3)+(in_buffer[2]<<6))+(0+(in_buffer[3]<<2)+(in_buffer[3]<<5))+(0-(in_buffer[4]<<0)-(in_buffer[4]<<2)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<1)+(in_buffer[5]<<4)+(in_buffer[5]<<5))-(0-(in_buffer[6]<<1)+(in_buffer[6]<<4))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<5)+(in_buffer[7]<<6))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<2))-(0-(in_buffer[9]<<0)+(in_buffer[9]<<4))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<3))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<6))-(0-(in_buffer[12]<<1)+(in_buffer[12]<<4))+(0+(in_buffer[13]<<1)+(in_buffer[13]<<4))+(0-(in_buffer[14]<<2)+(in_buffer[14]<<4)+(in_buffer[14]<<5))+(0+(in_buffer[15]<<1)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<4))+(0+(in_buffer[17]<<2))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<2)+(in_buffer[19]<<5))-(0-(in_buffer[20]<<2)+(in_buffer[20]<<5)+(in_buffer[20]<<6))-(0+(in_buffer[21]<<2)+(in_buffer[21]<<4))+(0-(in_buffer[22]<<3)+(in_buffer[22]<<6))-(0+(in_buffer[23]<<1)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<0));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight45;
assign in_buffer_weight45=0-(0+(in_buffer[0]<<1)+(in_buffer[0]<<2)+(in_buffer[0]<<6))-(0+(in_buffer[1]<<5))-(0-(in_buffer[2]<<1)+(in_buffer[2]<<3)+(in_buffer[2]<<4))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<2))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<5))+(0+(in_buffer[5]<<0))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<3))-(0+(in_buffer[7]<<0)-(in_buffer[7]<<2)+(in_buffer[7]<<6))+(0-(in_buffer[8]<<0)+(in_buffer[8]<<4)+(in_buffer[8]<<5))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<6))+(0+(in_buffer[10]<<2)+(in_buffer[10]<<5))+(0-(in_buffer[11]<<3)+(in_buffer[11]<<6))+(0-(in_buffer[12]<<1)-(in_buffer[12]<<3)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<5))-(0-(in_buffer[14]<<0)+(in_buffer[14]<<3)+(in_buffer[14]<<6))-(0+(in_buffer[15]<<0)-(in_buffer[15]<<3)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<5))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<3)+(in_buffer[17]<<5))-(0-(in_buffer[18]<<3)+(in_buffer[18]<<5)+(in_buffer[18]<<6))-(0+(in_buffer[19]<<0)+(in_buffer[19]<<2)-(in_buffer[19]<<4)+(in_buffer[19]<<7))-(0+(in_buffer[20]<<2)+(in_buffer[20]<<5))-(0-(in_buffer[21]<<0)+(in_buffer[21]<<4))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<1)+(in_buffer[22]<<4))+(0+(in_buffer[23]<<3)+(in_buffer[23]<<5)+(in_buffer[23]<<6))+(0+(in_buffer[24]<<2)+(in_buffer[24]<<4)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight46;
assign in_buffer_weight46=0+(0+(in_buffer[0]<<0)-(in_buffer[0]<<2)+(in_buffer[0]<<5)+(in_buffer[0]<<7))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<3)+(in_buffer[1]<<7))+(0-(in_buffer[2]<<0)-(in_buffer[2]<<3)+(in_buffer[2]<<7))-(0-(in_buffer[3]<<2)+(in_buffer[3]<<4)+(in_buffer[3]<<5))-(0-(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<3)+(in_buffer[4]<<6))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<3)+(in_buffer[5]<<5))-(0+(in_buffer[6]<<0))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<4)+(in_buffer[7]<<6))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<4)+(in_buffer[8]<<6))+(0-(in_buffer[9]<<0)-(in_buffer[9]<<2)+(in_buffer[9]<<5))-(0+(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<5))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<3)+(in_buffer[11]<<6))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<5))-(0+(in_buffer[13]<<1)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<2)+(in_buffer[14]<<4))-(0+(in_buffer[15]<<1)-(in_buffer[15]<<3)+(in_buffer[15]<<6))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<3))-(0+(in_buffer[17]<<2)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<3)+(in_buffer[18]<<4))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<3)+(in_buffer[19]<<5))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<3)+(in_buffer[20]<<5)+(in_buffer[20]<<6))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<5))+(0-(in_buffer[22]<<0)+(in_buffer[22]<<4))-(0+(in_buffer[23]<<2)+(in_buffer[23]<<4))-(0-(in_buffer[24]<<0)-(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight47;
assign in_buffer_weight47=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<4))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<4))-(0+(in_buffer[2]<<1)+(in_buffer[2]<<3))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<4))-(0+(in_buffer[4]<<0))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<4))+(0+(in_buffer[6]<<1))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<3))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<3))-(0-(in_buffer[9]<<0)+(in_buffer[9]<<4))-(0+(in_buffer[10]<<2))-(0-(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<4))-(0-(in_buffer[12]<<0)+(in_buffer[12]<<3))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2)+(in_buffer[13]<<4))-(0-(in_buffer[14]<<1)+(in_buffer[14]<<4))+(0+(in_buffer[15]<<1)+(in_buffer[15]<<2))-(0+(in_buffer[16]<<2)+(in_buffer[16]<<4))-(0+(in_buffer[17]<<2)+(in_buffer[17]<<3))+(0+(in_buffer[18]<<2))-(0+(in_buffer[19]<<3))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<4))-(0-(in_buffer[22]<<1)+(in_buffer[22]<<3)+(in_buffer[22]<<4))-(0-(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<1)+(in_buffer[24]<<4));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight48;
assign in_buffer_weight48=0+(0-(in_buffer[0]<<1)+(in_buffer[0]<<4)+(in_buffer[0]<<5))+(0-(in_buffer[2]<<0)+(in_buffer[2]<<4))+(0-(in_buffer[3]<<0)+(in_buffer[3]<<4))-(0-(in_buffer[4]<<1)+(in_buffer[4]<<5))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<5))+(0+(in_buffer[6]<<2)+(in_buffer[6]<<3))+(0-(in_buffer[7]<<1)+(in_buffer[7]<<4)+(in_buffer[7]<<5))+(0+(in_buffer[8]<<1)+(in_buffer[8]<<3))-(0+(in_buffer[9]<<5))+(0+(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<4)+(in_buffer[10]<<5))-(0+(in_buffer[11]<<1)+(in_buffer[11]<<5))-(0-(in_buffer[12]<<0)+(in_buffer[12]<<3))+(0+(in_buffer[13]<<2)+(in_buffer[13]<<4))+(0-(in_buffer[14]<<3)+(in_buffer[14]<<6))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<3))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<3)+(in_buffer[17]<<6))-(0-(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<6))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<5))-(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<5)+(in_buffer[22]<<6))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<2)+(in_buffer[23]<<6))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight49;
assign in_buffer_weight49=0-(0+(in_buffer[0]<<2)+(in_buffer[0]<<3)+(in_buffer[0]<<6))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<2))-(0+(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<5)+(in_buffer[2]<<6))-(0+(in_buffer[3]<<2))+(0-(in_buffer[4]<<1)+(in_buffer[4]<<4)+(in_buffer[4]<<5))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<6))+(0+(in_buffer[6]<<2)+(in_buffer[6]<<6))+(0+(in_buffer[7]<<3)+(in_buffer[7]<<4))+(0+(in_buffer[8]<<1)+(in_buffer[8]<<3)+(in_buffer[8]<<4))-(0-(in_buffer[9]<<1)+(in_buffer[9]<<6))+(0-(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<3))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3)+(in_buffer[11]<<6))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<5))-(0+(in_buffer[14]<<1))-(0+(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<5))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<6))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<5))-(0+(in_buffer[18]<<4))-(0+(in_buffer[19]<<3)+(in_buffer[19]<<4))-(0-(in_buffer[20]<<2)+(in_buffer[20]<<8))-(0+(in_buffer[21]<<3)+(in_buffer[21]<<5))+(0-(in_buffer[22]<<2)+(in_buffer[22]<<6))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)+(in_buffer[23]<<4)+(in_buffer[23]<<5))+(0+(in_buffer[24]<<2)+(in_buffer[24]<<3)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight50;
assign in_buffer_weight50=0+(0+(in_buffer[0]<<4)+(in_buffer[0]<<5))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<2)+(in_buffer[1]<<5))-(0-(in_buffer[2]<<0)+(in_buffer[2]<<5))+(0-(in_buffer[3]<<0)-(in_buffer[3]<<4)+(in_buffer[3]<<7))+(0+(in_buffer[4]<<0)-(in_buffer[4]<<3)+(in_buffer[4]<<5)+(in_buffer[4]<<6))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<5))-(0-(in_buffer[6]<<2)+(in_buffer[6]<<5)+(in_buffer[6]<<6))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<3)+(in_buffer[8]<<4))-(0+(in_buffer[9]<<1)+(in_buffer[9]<<5)+(in_buffer[9]<<7))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<1))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<2)+(in_buffer[11]<<5))+(0+(in_buffer[12]<<2)+(in_buffer[12]<<6))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<4))+(0+(in_buffer[14]<<1)+(in_buffer[14]<<3)+(in_buffer[14]<<4))+(0-(in_buffer[15]<<0)-(in_buffer[15]<<3)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<3)+(in_buffer[16]<<4))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<4))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<3))+(0-(in_buffer[19]<<0)-(in_buffer[19]<<2)-(in_buffer[19]<<4)+(in_buffer[19]<<7))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<2)+(in_buffer[20]<<5)+(in_buffer[20]<<6))-(0+(in_buffer[21]<<2)+(in_buffer[21]<<3))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<2)+(in_buffer[22]<<3))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<4))-(0-(in_buffer[24]<<1)+(in_buffer[24]<<4));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight51;
assign in_buffer_weight51=0+(0+(in_buffer[0]<<1)+(in_buffer[0]<<3)+(in_buffer[0]<<6))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<4)+(in_buffer[1]<<6))+(0-(in_buffer[2]<<0)+(in_buffer[2]<<5)+(in_buffer[2]<<6))+(0-(in_buffer[3]<<2)+(in_buffer[3]<<5)+(in_buffer[3]<<6))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<1)+(in_buffer[4]<<4))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<4))-(0+(in_buffer[6]<<1)+(in_buffer[6]<<6))-(0-(in_buffer[7]<<3)+(in_buffer[7]<<6))+(0+(in_buffer[8]<<6))+(0-(in_buffer[9]<<0)-(in_buffer[9]<<3)+(in_buffer[9]<<5)+(in_buffer[9]<<6))+(0+(in_buffer[10]<<1)+(in_buffer[10]<<3)+(in_buffer[10]<<4))-(0+(in_buffer[11]<<5))+(0+(in_buffer[12]<<3)+(in_buffer[12]<<4))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<1)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<5))+(0+(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<4)+(in_buffer[15]<<5))-(0-(in_buffer[16]<<1)+(in_buffer[16]<<5))+(0+(in_buffer[17]<<2)+(in_buffer[17]<<5))-(0-(in_buffer[18]<<2)+(in_buffer[18]<<5))-(0+(in_buffer[19]<<0)+(in_buffer[19]<<3)+(in_buffer[19]<<4))-(0+(in_buffer[20]<<2)+(in_buffer[20]<<3))+(0-(in_buffer[21]<<0)-(in_buffer[21]<<2)+(in_buffer[21]<<5))-(0+(in_buffer[22]<<2))+(0+(in_buffer[23]<<3)+(in_buffer[23]<<5))+(0-(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<4)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight52;
assign in_buffer_weight52=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3)+(in_buffer[0]<<7))-(0+(in_buffer[1]<<1)+(in_buffer[1]<<4)+(in_buffer[1]<<6))-(0-(in_buffer[2]<<0)+(in_buffer[2]<<3)+(in_buffer[2]<<4)+(in_buffer[2]<<7))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<7))-(0-(in_buffer[4]<<1)+(in_buffer[4]<<4)+(in_buffer[4]<<7))+(0+(in_buffer[5]<<4)+(in_buffer[5]<<5))+(0+(in_buffer[6]<<3)+(in_buffer[6]<<4))+(0-(in_buffer[7]<<0)+(in_buffer[7]<<4)+(in_buffer[7]<<5))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<1))+(0+(in_buffer[9]<<2)+(in_buffer[9]<<6))-(0+(in_buffer[10]<<4))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<1))+(0+(in_buffer[12]<<2)+(in_buffer[12]<<4))-(0+(in_buffer[13]<<1)+(in_buffer[13]<<2))-(0-(in_buffer[14]<<1)+(in_buffer[14]<<4))+(0+(in_buffer[15]<<3))+(0+(in_buffer[16]<<5))+(0+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<3))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<1)+(in_buffer[19]<<4))-(0+(in_buffer[20]<<3)+(in_buffer[20]<<7))-(0+(in_buffer[21]<<3)+(in_buffer[21]<<5))-(0-(in_buffer[22]<<1)-(in_buffer[22]<<3)+(in_buffer[22]<<5)+(in_buffer[22]<<6))-(0-(in_buffer[23]<<0)+(in_buffer[23]<<6))-(0-(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight53;
assign in_buffer_weight53=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<3))+(0-(in_buffer[1]<<3)+(in_buffer[1]<<6))+(0+(in_buffer[2]<<1)-(in_buffer[2]<<4)+(in_buffer[2]<<7))+(0-(in_buffer[3]<<1)+(in_buffer[3]<<4))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<4))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<5)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<3)+(in_buffer[6]<<5)+(in_buffer[6]<<6))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<4)+(in_buffer[7]<<6))+(0+(in_buffer[8]<<1)+(in_buffer[8]<<6))-(0-(in_buffer[9]<<0)-(in_buffer[9]<<2)+(in_buffer[9]<<4)+(in_buffer[9]<<5))-(0-(in_buffer[10]<<0)+(in_buffer[10]<<3))+(0+(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<5))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<5))+(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<1)+(in_buffer[14]<<3))-(0+(in_buffer[15]<<1)+(in_buffer[15]<<3))+(0+(in_buffer[16]<<2))+(0+(in_buffer[17]<<2))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<5))-(0+(in_buffer[19]<<1)+(in_buffer[19]<<3)+(in_buffer[19]<<4))+(0+(in_buffer[20]<<3))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<1))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<5))+(0+(in_buffer[23]<<2))+(0+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight54;
assign in_buffer_weight54=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<4))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<5))-(0-(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<6))-(0-(in_buffer[3]<<1)+(in_buffer[3]<<6))-(0+(in_buffer[4]<<6))+(0+(in_buffer[5]<<2)+(in_buffer[5]<<4)+(in_buffer[5]<<5))+(0+(in_buffer[6]<<1)+(in_buffer[6]<<3)+(in_buffer[6]<<5)+(in_buffer[6]<<6))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<5))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<3)+(in_buffer[8]<<4))+(0-(in_buffer[9]<<1)+(in_buffer[9]<<3)+(in_buffer[9]<<4))-(0+(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<6))+(0+(in_buffer[12]<<1)+(in_buffer[12]<<3))-(0+(in_buffer[13]<<0))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<1)+(in_buffer[14]<<5))-(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<4)+(in_buffer[15]<<5))-(0+(in_buffer[16]<<1))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<3)+(in_buffer[17]<<6))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<3)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<2))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<3)+(in_buffer[20]<<4))+(0-(in_buffer[21]<<1)+(in_buffer[21]<<4))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<3))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)+(in_buffer[23]<<4)+(in_buffer[23]<<5))-(0+(in_buffer[24]<<1));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight55;
assign in_buffer_weight55=0-(0+(in_buffer[0]<<2)+(in_buffer[0]<<6))-(0+(in_buffer[2]<<2)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<5)+(in_buffer[3]<<6))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<3)-(in_buffer[4]<<5)+(in_buffer[4]<<8))+(0+(in_buffer[5]<<0)+(in_buffer[5]<<1)+(in_buffer[5]<<4)+(in_buffer[5]<<5))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<4))+(0-(in_buffer[7]<<1)+(in_buffer[7]<<3)+(in_buffer[7]<<4))+(0+(in_buffer[8]<<1)+(in_buffer[8]<<3)+(in_buffer[8]<<6))-(0+(in_buffer[9]<<1)+(in_buffer[9]<<4))+(0-(in_buffer[10]<<0)+(in_buffer[10]<<4))-(0+(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<6))-(0-(in_buffer[12]<<0)+(in_buffer[12]<<5))+(0+(in_buffer[13]<<3))+(0+(in_buffer[14]<<1)+(in_buffer[14]<<3)+(in_buffer[14]<<4))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<3))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<3))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<4))-(0+(in_buffer[19]<<4))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<4)+(in_buffer[20]<<5))+(0-(in_buffer[21]<<2)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<2))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<3)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<5)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight56;
assign in_buffer_weight56=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<5))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<4))-(0-(in_buffer[2]<<0)+(in_buffer[2]<<3)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<5))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<1))+(0+(in_buffer[5]<<0)+(in_buffer[5]<<1)+(in_buffer[5]<<4))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<4))+(0-(in_buffer[7]<<2)+(in_buffer[7]<<6))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<2)+(in_buffer[8]<<3)+(in_buffer[8]<<6))+(0+(in_buffer[9]<<4)+(in_buffer[9]<<5))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<3))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<5))-(0+(in_buffer[12]<<1)+(in_buffer[12]<<5))-(0-(in_buffer[13]<<1)+(in_buffer[13]<<4)+(in_buffer[13]<<6))+(0+(in_buffer[14]<<1)+(in_buffer[14]<<3)+(in_buffer[14]<<4))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3)+(in_buffer[15]<<5))+(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<5))-(0-(in_buffer[17]<<0)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<3))+(0+(in_buffer[19]<<1)-(in_buffer[19]<<3)+(in_buffer[19]<<6))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<3)+(in_buffer[20]<<5))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<5))+(0-(in_buffer[22]<<0)+(in_buffer[22]<<2)+(in_buffer[22]<<3))+(0+(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<5))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<2));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight57;
assign in_buffer_weight57=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<5))-(0-(in_buffer[2]<<1)+(in_buffer[2]<<5)+(in_buffer[2]<<6))+(0+(in_buffer[3]<<2)+(in_buffer[3]<<4)+(in_buffer[3]<<6))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<2)+(in_buffer[4]<<6))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3))+(0-(in_buffer[6]<<1)+(in_buffer[6]<<4)+(in_buffer[6]<<5))+(0-(in_buffer[7]<<1)+(in_buffer[7]<<5))+(0-(in_buffer[8]<<0)+(in_buffer[8]<<5))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<3)+(in_buffer[9]<<5))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<3)+(in_buffer[10]<<4))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<3))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<1)+(in_buffer[12]<<6))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<6))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<4)+(in_buffer[14]<<7))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<4))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<4))+(0+(in_buffer[18]<<2)+(in_buffer[18]<<3))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<6))+(0+(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<1)+(in_buffer[21]<<4))+(0-(in_buffer[22]<<2)+(in_buffer[22]<<5))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<4))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight58;
assign in_buffer_weight58=0+(0+(in_buffer[0]<<4)+(in_buffer[0]<<6)+(in_buffer[0]<<7))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<2)+(in_buffer[1]<<7))-(0+(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<4))+(0+(in_buffer[4]<<2)+(in_buffer[4]<<3))-(0+(in_buffer[5]<<3)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<3)+(in_buffer[6]<<5)+(in_buffer[6]<<6))-(0-(in_buffer[7]<<1)+(in_buffer[7]<<3)+(in_buffer[7]<<4))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<2))-(0-(in_buffer[9]<<0)+(in_buffer[9]<<3)+(in_buffer[9]<<6))+(0-(in_buffer[10]<<1)+(in_buffer[10]<<4))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3)+(in_buffer[11]<<6))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<3)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<1)+(in_buffer[14]<<2)+(in_buffer[14]<<5))+(0+(in_buffer[15]<<4)+(in_buffer[15]<<5))+(0+(in_buffer[16]<<1))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<1))+(0+(in_buffer[18]<<3)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<1))-(0+(in_buffer[20]<<2)+(in_buffer[20]<<4)+(in_buffer[20]<<5))-(0+(in_buffer[21]<<1))-(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<4)+(in_buffer[23]<<5))-(0-(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<7));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight59;
assign in_buffer_weight59=0+(0+(in_buffer[1]<<1)+(in_buffer[1]<<2))-(0+(in_buffer[2]<<1))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<3)+(in_buffer[3]<<4))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<1)+(in_buffer[4]<<4))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<4))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<4))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<2))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<2))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<3))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<3))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<1))-(0+(in_buffer[12]<<3))+(0+(in_buffer[13]<<0)+(in_buffer[13]<<2))-(0-(in_buffer[14]<<0)+(in_buffer[14]<<3)+(in_buffer[14]<<4))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<4))-(0+(in_buffer[16]<<3))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4))+(0-(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<3))-(0-(in_buffer[19]<<1)+(in_buffer[19]<<4))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2))-(0+(in_buffer[21]<<1)+(in_buffer[21]<<2))+(0+(in_buffer[22]<<3))+(0-(in_buffer[23]<<0)+(in_buffer[23]<<3))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight60;
assign in_buffer_weight60=0-(0+(in_buffer[0]<<0)-(in_buffer[0]<<5)+(in_buffer[0]<<8))-(0+(in_buffer[1]<<1)-(in_buffer[1]<<3)+(in_buffer[1]<<5)+(in_buffer[1]<<6))+(0+(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<2)+(in_buffer[3]<<3))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<3)+(in_buffer[4]<<6))+(0+(in_buffer[5]<<2)-(in_buffer[5]<<4)+(in_buffer[5]<<7))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<4)+(in_buffer[6]<<5))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<3))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<2))+(0+(in_buffer[9]<<3)+(in_buffer[9]<<6))+(0+(in_buffer[10]<<1)+(in_buffer[10]<<3))-(0-(in_buffer[11]<<2)+(in_buffer[11]<<5))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<3)+(in_buffer[12]<<5))+(0-(in_buffer[13]<<2)+(in_buffer[13]<<4)+(in_buffer[13]<<5))-(0-(in_buffer[14]<<0)+(in_buffer[14]<<4)+(in_buffer[14]<<5))-(0+(in_buffer[15]<<3)+(in_buffer[15]<<5))-(0-(in_buffer[16]<<2)+(in_buffer[16]<<4)+(in_buffer[16]<<5))-(0-(in_buffer[17]<<1)+(in_buffer[17]<<4))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<5))-(0+(in_buffer[19]<<0)-(in_buffer[19]<<3)+(in_buffer[19]<<5)+(in_buffer[19]<<6))-(0+(in_buffer[20]<<3))+(0-(in_buffer[21]<<1)+(in_buffer[21]<<4))+(0-(in_buffer[22]<<1)+(in_buffer[22]<<3)+(in_buffer[22]<<4))+(0+(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<5))+(0-(in_buffer[24]<<2)+(in_buffer[24]<<5)+(in_buffer[24]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight61;
assign in_buffer_weight61=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<5))+(0+(in_buffer[1]<<4))-(0+(in_buffer[2]<<4)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<3))+(0+(in_buffer[4]<<3))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<2))-(0-(in_buffer[6]<<2)+(in_buffer[6]<<4)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<1)+(in_buffer[7]<<4))+(0-(in_buffer[8]<<3)+(in_buffer[8]<<5)+(in_buffer[8]<<6))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<3))-(0+(in_buffer[10]<<4))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<4))+(0+(in_buffer[12]<<4)+(in_buffer[12]<<5))+(0+(in_buffer[13]<<2)+(in_buffer[13]<<4)+(in_buffer[13]<<5))+(0-(in_buffer[14]<<3)+(in_buffer[14]<<6))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<4)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<1)+(in_buffer[17]<<3)+(in_buffer[17]<<4))-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<6))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<2))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<3)+(in_buffer[20]<<6))+(0+(in_buffer[22]<<3)+(in_buffer[22]<<5))-(0-(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<3)+(in_buffer[23]<<6))-(0+(in_buffer[24]<<2)+(in_buffer[24]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight62;
assign in_buffer_weight62=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<7))-(0-(in_buffer[1]<<0)+(in_buffer[1]<<3))+(0-(in_buffer[2]<<2)+(in_buffer[2]<<4)+(in_buffer[2]<<5))-(0+(in_buffer[3]<<0)-(in_buffer[3]<<3)+(in_buffer[3]<<7))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<4))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3)+(in_buffer[5]<<6))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<3)+(in_buffer[6]<<5))+(0+(in_buffer[7]<<1))+(0+(in_buffer[9]<<0)-(in_buffer[9]<<3)+(in_buffer[9]<<6))-(0+(in_buffer[10]<<2)+(in_buffer[10]<<4)+(in_buffer[10]<<5))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<4)+(in_buffer[11]<<5))-(0+(in_buffer[12]<<1))+(0+(in_buffer[13]<<3)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<2)+(in_buffer[14]<<3)+(in_buffer[14]<<6))+(0+(in_buffer[15]<<2))+(0-(in_buffer[16]<<0)-(in_buffer[16]<<2)+(in_buffer[16]<<4)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<5))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<2)+(in_buffer[18]<<5))-(0+(in_buffer[19]<<0)-(in_buffer[19]<<2)+(in_buffer[19]<<6))+(0+(in_buffer[20]<<1))+(0+(in_buffer[21]<<1))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<3))-(0+(in_buffer[23]<<2)+(in_buffer[23]<<3))+(0+(in_buffer[24]<<0)-(in_buffer[24]<<2)+(in_buffer[24]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight63;
assign in_buffer_weight63=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<4)+(in_buffer[0]<<7))-(0-(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<3)+(in_buffer[1]<<7))+(0-(in_buffer[2]<<1)+(in_buffer[2]<<4)+(in_buffer[2]<<5))-(0-(in_buffer[3]<<3)+(in_buffer[3]<<6))-(0+(in_buffer[4]<<2)-(in_buffer[4]<<4)+(in_buffer[4]<<7))+(0+(in_buffer[5]<<3)+(in_buffer[5]<<5))+(0-(in_buffer[6]<<1)+(in_buffer[6]<<3)+(in_buffer[6]<<4))+(0+(in_buffer[7]<<2)+(in_buffer[7]<<3))+(0+(in_buffer[8]<<2)+(in_buffer[8]<<6))+(0-(in_buffer[9]<<0)+(in_buffer[9]<<5))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<3)+(in_buffer[10]<<5)+(in_buffer[10]<<6))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<3))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<1)+(in_buffer[13]<<6))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<4)+(in_buffer[14]<<5))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<1))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4)+(in_buffer[17]<<5))+(0-(in_buffer[18]<<0)+(in_buffer[18]<<3)+(in_buffer[18]<<5)+(in_buffer[18]<<6))-(0-(in_buffer[19]<<0)-(in_buffer[19]<<3)+(in_buffer[19]<<6))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<3)+(in_buffer[20]<<7))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<4))+(0-(in_buffer[22]<<3)+(in_buffer[22]<<6))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<4)+(in_buffer[23]<<6))-(0-(in_buffer[24]<<1)-(in_buffer[24]<<3)-(in_buffer[24]<<5)+(in_buffer[24]<<7)+(in_buffer[24]<<8));
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
wire signed [DATA_WIDTH-1:0]   weight_bias10;
wire signed [DATA_WIDTH-1:0]   weight_bias11;
wire signed [DATA_WIDTH-1:0]   weight_bias12;
wire signed [DATA_WIDTH-1:0]   weight_bias13;
wire signed [DATA_WIDTH-1:0]   weight_bias14;
wire signed [DATA_WIDTH-1:0]   weight_bias15;
wire signed [DATA_WIDTH-1:0]   weight_bias16;
wire signed [DATA_WIDTH-1:0]   weight_bias17;
wire signed [DATA_WIDTH-1:0]   weight_bias18;
wire signed [DATA_WIDTH-1:0]   weight_bias19;
wire signed [DATA_WIDTH-1:0]   weight_bias20;
wire signed [DATA_WIDTH-1:0]   weight_bias21;
wire signed [DATA_WIDTH-1:0]   weight_bias22;
wire signed [DATA_WIDTH-1:0]   weight_bias23;
wire signed [DATA_WIDTH-1:0]   weight_bias24;
wire signed [DATA_WIDTH-1:0]   weight_bias25;
wire signed [DATA_WIDTH-1:0]   weight_bias26;
wire signed [DATA_WIDTH-1:0]   weight_bias27;
wire signed [DATA_WIDTH-1:0]   weight_bias28;
wire signed [DATA_WIDTH-1:0]   weight_bias29;
wire signed [DATA_WIDTH-1:0]   weight_bias30;
wire signed [DATA_WIDTH-1:0]   weight_bias31;
wire signed [DATA_WIDTH-1:0]   weight_bias32;
wire signed [DATA_WIDTH-1:0]   weight_bias33;
wire signed [DATA_WIDTH-1:0]   weight_bias34;
wire signed [DATA_WIDTH-1:0]   weight_bias35;
wire signed [DATA_WIDTH-1:0]   weight_bias36;
wire signed [DATA_WIDTH-1:0]   weight_bias37;
wire signed [DATA_WIDTH-1:0]   weight_bias38;
wire signed [DATA_WIDTH-1:0]   weight_bias39;
wire signed [DATA_WIDTH-1:0]   weight_bias40;
wire signed [DATA_WIDTH-1:0]   weight_bias41;
wire signed [DATA_WIDTH-1:0]   weight_bias42;
wire signed [DATA_WIDTH-1:0]   weight_bias43;
wire signed [DATA_WIDTH-1:0]   weight_bias44;
wire signed [DATA_WIDTH-1:0]   weight_bias45;
wire signed [DATA_WIDTH-1:0]   weight_bias46;
wire signed [DATA_WIDTH-1:0]   weight_bias47;
wire signed [DATA_WIDTH-1:0]   weight_bias48;
wire signed [DATA_WIDTH-1:0]   weight_bias49;
wire signed [DATA_WIDTH-1:0]   weight_bias50;
wire signed [DATA_WIDTH-1:0]   weight_bias51;
wire signed [DATA_WIDTH-1:0]   weight_bias52;
wire signed [DATA_WIDTH-1:0]   weight_bias53;
wire signed [DATA_WIDTH-1:0]   weight_bias54;
wire signed [DATA_WIDTH-1:0]   weight_bias55;
wire signed [DATA_WIDTH-1:0]   weight_bias56;
wire signed [DATA_WIDTH-1:0]   weight_bias57;
wire signed [DATA_WIDTH-1:0]   weight_bias58;
wire signed [DATA_WIDTH-1:0]   weight_bias59;
wire signed [DATA_WIDTH-1:0]   weight_bias60;
wire signed [DATA_WIDTH-1:0]   weight_bias61;
wire signed [DATA_WIDTH-1:0]   weight_bias62;
wire signed [DATA_WIDTH-1:0]   weight_bias63;
assign weight_bias0=in_buffer_weight0+(0);
assign weight_bias1=in_buffer_weight1+(39);
assign weight_bias2=in_buffer_weight2+(26);
assign weight_bias3=in_buffer_weight3+(-27);
assign weight_bias4=in_buffer_weight4+(2);
assign weight_bias5=in_buffer_weight5+(7);
assign weight_bias6=in_buffer_weight6+(-26);
assign weight_bias7=in_buffer_weight7+(-20);
assign weight_bias8=in_buffer_weight8+(-15);
assign weight_bias9=in_buffer_weight9+(27);
assign weight_bias10=in_buffer_weight10+(-6);
assign weight_bias11=in_buffer_weight11+(-5);
assign weight_bias12=in_buffer_weight12+(108);
assign weight_bias13=in_buffer_weight13+(-21);
assign weight_bias14=in_buffer_weight14+(16);
assign weight_bias15=in_buffer_weight15+(-3);
assign weight_bias16=in_buffer_weight16+(210);
assign weight_bias17=in_buffer_weight17+(54);
assign weight_bias18=in_buffer_weight18+(61);
assign weight_bias19=in_buffer_weight19+(12);
assign weight_bias20=in_buffer_weight20+(8);
assign weight_bias21=in_buffer_weight21+(44);
assign weight_bias22=in_buffer_weight22+(10);
assign weight_bias23=in_buffer_weight23+(47);
assign weight_bias24=in_buffer_weight24+(-32);
assign weight_bias25=in_buffer_weight25+(-31);
assign weight_bias26=in_buffer_weight26+(-22);
assign weight_bias27=in_buffer_weight27+(41);
assign weight_bias28=in_buffer_weight28+(-72);
assign weight_bias29=in_buffer_weight29+(-48);
assign weight_bias30=in_buffer_weight30+(-99);
assign weight_bias31=in_buffer_weight31+(5);
assign weight_bias32=in_buffer_weight32+(-2);
assign weight_bias33=in_buffer_weight33+(55);
assign weight_bias34=in_buffer_weight34+(81);
assign weight_bias35=in_buffer_weight35+(36);
assign weight_bias36=in_buffer_weight36+(-55);
assign weight_bias37=in_buffer_weight37+(6);
assign weight_bias38=in_buffer_weight38+(57);
assign weight_bias39=in_buffer_weight39+(13);
assign weight_bias40=in_buffer_weight40+(-17);
assign weight_bias41=in_buffer_weight41+(-35);
assign weight_bias42=in_buffer_weight42+(50);
assign weight_bias43=in_buffer_weight43+(-31);
assign weight_bias44=in_buffer_weight44+(29);
assign weight_bias45=in_buffer_weight45+(26);
assign weight_bias46=in_buffer_weight46+(-71);
assign weight_bias47=in_buffer_weight47+(-24);
assign weight_bias48=in_buffer_weight48+(50);
assign weight_bias49=in_buffer_weight49+(34);
assign weight_bias50=in_buffer_weight50+(55);
assign weight_bias51=in_buffer_weight51+(-19);
assign weight_bias52=in_buffer_weight52+(115);
assign weight_bias53=in_buffer_weight53+(-77);
assign weight_bias54=in_buffer_weight54+(66);
assign weight_bias55=in_buffer_weight55+(30);
assign weight_bias56=in_buffer_weight56+(-33);
assign weight_bias57=in_buffer_weight57+(10);
assign weight_bias58=in_buffer_weight58+(3);
assign weight_bias59=in_buffer_weight59+(-6);
assign weight_bias60=in_buffer_weight60+(6);
assign weight_bias61=in_buffer_weight61+(-19);
assign weight_bias62=in_buffer_weight62+(66);
assign weight_bias63=in_buffer_weight63+(52);
wire signed [DATA_WIDTH-1:0]   bias_relu0;
wire signed [DATA_WIDTH-1:0]   bias_relu1;
wire signed [DATA_WIDTH-1:0]   bias_relu2;
wire signed [DATA_WIDTH-1:0]   bias_relu3;
wire signed [DATA_WIDTH-1:0]   bias_relu4;
wire signed [DATA_WIDTH-1:0]   bias_relu5;
wire signed [DATA_WIDTH-1:0]   bias_relu6;
wire signed [DATA_WIDTH-1:0]   bias_relu7;
wire signed [DATA_WIDTH-1:0]   bias_relu8;
wire signed [DATA_WIDTH-1:0]   bias_relu9;
wire signed [DATA_WIDTH-1:0]   bias_relu10;
wire signed [DATA_WIDTH-1:0]   bias_relu11;
wire signed [DATA_WIDTH-1:0]   bias_relu12;
wire signed [DATA_WIDTH-1:0]   bias_relu13;
wire signed [DATA_WIDTH-1:0]   bias_relu14;
wire signed [DATA_WIDTH-1:0]   bias_relu15;
wire signed [DATA_WIDTH-1:0]   bias_relu16;
wire signed [DATA_WIDTH-1:0]   bias_relu17;
wire signed [DATA_WIDTH-1:0]   bias_relu18;
wire signed [DATA_WIDTH-1:0]   bias_relu19;
wire signed [DATA_WIDTH-1:0]   bias_relu20;
wire signed [DATA_WIDTH-1:0]   bias_relu21;
wire signed [DATA_WIDTH-1:0]   bias_relu22;
wire signed [DATA_WIDTH-1:0]   bias_relu23;
wire signed [DATA_WIDTH-1:0]   bias_relu24;
wire signed [DATA_WIDTH-1:0]   bias_relu25;
wire signed [DATA_WIDTH-1:0]   bias_relu26;
wire signed [DATA_WIDTH-1:0]   bias_relu27;
wire signed [DATA_WIDTH-1:0]   bias_relu28;
wire signed [DATA_WIDTH-1:0]   bias_relu29;
wire signed [DATA_WIDTH-1:0]   bias_relu30;
wire signed [DATA_WIDTH-1:0]   bias_relu31;
wire signed [DATA_WIDTH-1:0]   bias_relu32;
wire signed [DATA_WIDTH-1:0]   bias_relu33;
wire signed [DATA_WIDTH-1:0]   bias_relu34;
wire signed [DATA_WIDTH-1:0]   bias_relu35;
wire signed [DATA_WIDTH-1:0]   bias_relu36;
wire signed [DATA_WIDTH-1:0]   bias_relu37;
wire signed [DATA_WIDTH-1:0]   bias_relu38;
wire signed [DATA_WIDTH-1:0]   bias_relu39;
wire signed [DATA_WIDTH-1:0]   bias_relu40;
wire signed [DATA_WIDTH-1:0]   bias_relu41;
wire signed [DATA_WIDTH-1:0]   bias_relu42;
wire signed [DATA_WIDTH-1:0]   bias_relu43;
wire signed [DATA_WIDTH-1:0]   bias_relu44;
wire signed [DATA_WIDTH-1:0]   bias_relu45;
wire signed [DATA_WIDTH-1:0]   bias_relu46;
wire signed [DATA_WIDTH-1:0]   bias_relu47;
wire signed [DATA_WIDTH-1:0]   bias_relu48;
wire signed [DATA_WIDTH-1:0]   bias_relu49;
wire signed [DATA_WIDTH-1:0]   bias_relu50;
wire signed [DATA_WIDTH-1:0]   bias_relu51;
wire signed [DATA_WIDTH-1:0]   bias_relu52;
wire signed [DATA_WIDTH-1:0]   bias_relu53;
wire signed [DATA_WIDTH-1:0]   bias_relu54;
wire signed [DATA_WIDTH-1:0]   bias_relu55;
wire signed [DATA_WIDTH-1:0]   bias_relu56;
wire signed [DATA_WIDTH-1:0]   bias_relu57;
wire signed [DATA_WIDTH-1:0]   bias_relu58;
wire signed [DATA_WIDTH-1:0]   bias_relu59;
wire signed [DATA_WIDTH-1:0]   bias_relu60;
wire signed [DATA_WIDTH-1:0]   bias_relu61;
wire signed [DATA_WIDTH-1:0]   bias_relu62;
wire signed [DATA_WIDTH-1:0]   bias_relu63;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign bias_relu32=(weight_bias32[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias32;
assign bias_relu33=(weight_bias33[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias33;
assign bias_relu34=(weight_bias34[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias34;
assign bias_relu35=(weight_bias35[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias35;
assign bias_relu36=(weight_bias36[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias36;
assign bias_relu37=(weight_bias37[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias37;
assign bias_relu38=(weight_bias38[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias38;
assign bias_relu39=(weight_bias39[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias39;
assign bias_relu40=(weight_bias40[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias40;
assign bias_relu41=(weight_bias41[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias41;
assign bias_relu42=(weight_bias42[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias42;
assign bias_relu43=(weight_bias43[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias43;
assign bias_relu44=(weight_bias44[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias44;
assign bias_relu45=(weight_bias45[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias45;
assign bias_relu46=(weight_bias46[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias46;
assign bias_relu47=(weight_bias47[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias47;
assign bias_relu48=(weight_bias48[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias48;
assign bias_relu49=(weight_bias49[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias49;
assign bias_relu50=(weight_bias50[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias50;
assign bias_relu51=(weight_bias51[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias51;
assign bias_relu52=(weight_bias52[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias52;
assign bias_relu53=(weight_bias53[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias53;
assign bias_relu54=(weight_bias54[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias54;
assign bias_relu55=(weight_bias55[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias55;
assign bias_relu56=(weight_bias56[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias56;
assign bias_relu57=(weight_bias57[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias57;
assign bias_relu58=(weight_bias58[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias58;
assign bias_relu59=(weight_bias59[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias59;
assign bias_relu60=(weight_bias60[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias60;
assign bias_relu61=(weight_bias61[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias61;
assign bias_relu62=(weight_bias62[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias62;
assign bias_relu63=(weight_bias63[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias63;
assign layer_out={bias_relu63,bias_relu62,bias_relu61,bias_relu60,bias_relu59,bias_relu58,bias_relu57,bias_relu56,bias_relu55,bias_relu54,bias_relu53,bias_relu52,bias_relu51,bias_relu50,bias_relu49,bias_relu48,bias_relu47,bias_relu46,bias_relu45,bias_relu44,bias_relu43,bias_relu42,bias_relu41,bias_relu40,bias_relu39,bias_relu38,bias_relu37,bias_relu36,bias_relu35,bias_relu34,bias_relu33,bias_relu32,bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule