`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/22/2022 01:25:54 PM
// Design Name: 
// Module Name: n13sys4x4_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module n13sys4x4_testbench(

    );
    
    reg [5:0] word0,word1,word2,word3,word4,word5,word6,word7,word8,word9,word10,word11,word12,word13,word14,word15;
    wire [2:0]d_word0,d_word1,d_word2,d_word3,d_word4,d_word5,d_word6,d_word7,d_word8,d_word9,d_word10,d_word11,d_word12,d_word13,d_word14,d_word15;
    n13sys_4x4 DUT_n13(.IN0(word0),.IN1(word1),.IN2(word2),.IN3(word3),.IN4(word4),.IN5(word5),.IN6(word6),.IN7(word7),.IN8(word8),.IN9(word9),.IN10(word10),.IN11(word11),.IN12(word12),.IN13(word13),.IN14(word14),.IN15(word15),.OUT0(d_word0),.OUT1(d_word1),.OUT2(d_word2),.OUT3(d_word3),.OUT4(d_word4),.OUT5(d_word5),.OUT6(d_word6),.OUT7(d_word7),.OUT8(d_word8),.OUT9(d_word9),.OUT10(d_word10),.OUT11(d_word11),.OUT12(d_word12),.OUT13(d_word13),.OUT14(d_word14),.OUT15(d_word15));
    
    initial begin 
    
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
	#10 word0='d13;
	 #10 word0='d26;
	 #10 word0='d39;
	 #10 word0='d52;
    #10 word0='d1;
    #10 word0='d12;
    #10 word0='d27;
    #10 word0='d38;
    #10 word0='d53;
    #10 word0='d2;
    #10 word0='d15;
    #10 word0='d24;
    #10 word0='d37;
    #10 word0='d54;
    #10 word0='d4;
    #10 word0='d9;
    #10 word0='d30;
    #10 word0='d35;
    #10 word0='d48;
    #10 word0='d8;
    #10 word0='d5;
    #10 word0='d18;
    #10 word0='d47;
    #10 word0='d60;
    #10 word0='d16;
    #10 word0='d29;
    #10 word0='d10;
    #10 word0='d55;
    #10 word0='d36;
    #10 word0='d32;
    #10 word0='d45;
    #10 word0='d58;
    #10 word0='d7;
    #10 word0='d20;

/*
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word0='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word1='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word2='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word3='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word4='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word5='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word6='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word7='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word8='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word9='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word10='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word11='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word12='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word13='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word14='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
#10 word15='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;
*/
    
//word1
#20 $stop;
    end
endmodule
