module layer0_cnn_144_25x64x10
(
    input clk,
    input rst,
    input [475-1:0] layer_in,
    input valid,
    output  reg ready,
    output [27*64-1:0] layer_out
);
parameter DATA_WIDTH = 27;
parameter INPUT_DATA_CNT   =   25;
reg    signed [DATA_WIDTH-1:0]  in_buffer[0:INPUT_DATA_CNT-1];
genvar j;
generate
for(j=0;j<INPUT_DATA_CNT;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=layer_in[j*19+18:j*19+0];
                    end
            end
    end
endgenerate
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=$signed(in_buffer[0]*(9))+$signed(in_buffer[1]*(21))+$signed(in_buffer[2]*(6))+$signed(in_buffer[3]*(5))+$signed(in_buffer[4]*(-52))+$signed(in_buffer[5]*(3))+$signed(in_buffer[6]*(-3))+$signed(in_buffer[7]*(4))+$signed(in_buffer[8]*(8))+$signed(in_buffer[9]*(-9))+$signed(in_buffer[10]*(-7))+$signed(in_buffer[11]*(-106))+$signed(in_buffer[12]*(-85))+$signed(in_buffer[13]*(4))+$signed(in_buffer[14]*(45))+$signed(in_buffer[15]*(38))+$signed(in_buffer[16]*(-3))+$signed(in_buffer[17]*(45))+$signed(in_buffer[18]*(82))+$signed(in_buffer[19]*(19))+$signed(in_buffer[20]*(15))+$signed(in_buffer[21]*(60))+$signed(in_buffer[22]*(5))+$signed(in_buffer[23]*(-6))+$signed(in_buffer[24]*(-28));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=$signed(in_buffer[0]*(33))+$signed(in_buffer[1]*(125))+$signed(in_buffer[2]*(100))+$signed(in_buffer[3]*(22))+$signed(in_buffer[4]*(-40))+$signed(in_buffer[5]*(38))+$signed(in_buffer[6]*(16))+$signed(in_buffer[7]*(-15))+$signed(in_buffer[8]*(-38))+$signed(in_buffer[9]*(-67))+$signed(in_buffer[10]*(-86))+$signed(in_buffer[11]*(-27))+$signed(in_buffer[12]*(-13))+$signed(in_buffer[13]*(-30))+$signed(in_buffer[14]*(29))+$signed(in_buffer[15]*(-56))+$signed(in_buffer[16]*(-61))+$signed(in_buffer[17]*(-13))+$signed(in_buffer[18]*(24))+$signed(in_buffer[19]*(41))+$signed(in_buffer[20]*(112))+$signed(in_buffer[21]*(65))+$signed(in_buffer[22]*(31))+$signed(in_buffer[23]*(58))+$signed(in_buffer[24]*(43));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=$signed(in_buffer[0]*(-24))+$signed(in_buffer[1]*(-49))+$signed(in_buffer[2]*(-59))+$signed(in_buffer[3]*(-47))+$signed(in_buffer[4]*(29))+$signed(in_buffer[5]*(-2))+$signed(in_buffer[6]*(31))+$signed(in_buffer[7]*(56))+$signed(in_buffer[8]*(-38))+$signed(in_buffer[9]*(3))+$signed(in_buffer[10]*(-32))+$signed(in_buffer[11]*(-13))+$signed(in_buffer[12]*(-3))+$signed(in_buffer[13]*(58))+$signed(in_buffer[14]*(34))+$signed(in_buffer[15]*(6))+$signed(in_buffer[16]*(-5))+$signed(in_buffer[17]*(-23))+$signed(in_buffer[18]*(18))+$signed(in_buffer[19]*(1))+$signed(in_buffer[20]*(54))+$signed(in_buffer[21]*(-4))+$signed(in_buffer[22]*(0))+$signed(in_buffer[23]*(34))+$signed(in_buffer[24]*(39));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=$signed(in_buffer[0]*(9))+$signed(in_buffer[1]*(4))+$signed(in_buffer[2]*(13))+$signed(in_buffer[3]*(-15))+$signed(in_buffer[4]*(12))+$signed(in_buffer[5]*(36))+$signed(in_buffer[6]*(-16))+$signed(in_buffer[7]*(27))+$signed(in_buffer[8]*(23))+$signed(in_buffer[9]*(53))+$signed(in_buffer[10]*(42))+$signed(in_buffer[11]*(1))+$signed(in_buffer[12]*(-26))+$signed(in_buffer[13]*(-40))+$signed(in_buffer[14]*(114))+$signed(in_buffer[15]*(20))+$signed(in_buffer[16]*(-6))+$signed(in_buffer[17]*(-67))+$signed(in_buffer[18]*(44))+$signed(in_buffer[19]*(-22))+$signed(in_buffer[20]*(-32))+$signed(in_buffer[21]*(-9))+$signed(in_buffer[22]*(55))+$signed(in_buffer[23]*(48))+$signed(in_buffer[24]*(-27));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=$signed(in_buffer[0]*(7))+$signed(in_buffer[1]*(-33))+$signed(in_buffer[2]*(-72))+$signed(in_buffer[3]*(-31))+$signed(in_buffer[4]*(21))+$signed(in_buffer[5]*(-19))+$signed(in_buffer[6]*(1))+$signed(in_buffer[7]*(14))+$signed(in_buffer[8]*(47))+$signed(in_buffer[9]*(-52))+$signed(in_buffer[10]*(61))+$signed(in_buffer[11]*(19))+$signed(in_buffer[12]*(-38))+$signed(in_buffer[13]*(56))+$signed(in_buffer[14]*(15))+$signed(in_buffer[15]*(7))+$signed(in_buffer[16]*(-2))+$signed(in_buffer[17]*(23))+$signed(in_buffer[18]*(18))+$signed(in_buffer[19]*(-11))+$signed(in_buffer[20]*(-61))+$signed(in_buffer[21]*(45))+$signed(in_buffer[22]*(-24))+$signed(in_buffer[23]*(-66))+$signed(in_buffer[24]*(-147));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=$signed(in_buffer[0]*(-32))+$signed(in_buffer[1]*(-12))+$signed(in_buffer[2]*(28))+$signed(in_buffer[3]*(67))+$signed(in_buffer[4]*(21))+$signed(in_buffer[5]*(-15))+$signed(in_buffer[6]*(7))+$signed(in_buffer[7]*(-18))+$signed(in_buffer[8]*(-12))+$signed(in_buffer[9]*(68))+$signed(in_buffer[10]*(-12))+$signed(in_buffer[11]*(-8))+$signed(in_buffer[12]*(-101))+$signed(in_buffer[13]*(36))+$signed(in_buffer[14]*(46))+$signed(in_buffer[15]*(-40))+$signed(in_buffer[16]*(-1))+$signed(in_buffer[17]*(-11))+$signed(in_buffer[18]*(-14))+$signed(in_buffer[19]*(-28))+$signed(in_buffer[20]*(3))+$signed(in_buffer[21]*(96))+$signed(in_buffer[22]*(-20))+$signed(in_buffer[23]*(-45))+$signed(in_buffer[24]*(-5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=$signed(in_buffer[0]*(-13))+$signed(in_buffer[1]*(-92))+$signed(in_buffer[2]*(-9))+$signed(in_buffer[3]*(0))+$signed(in_buffer[4]*(0))+$signed(in_buffer[5]*(15))+$signed(in_buffer[6]*(-48))+$signed(in_buffer[7]*(47))+$signed(in_buffer[8]*(-5))+$signed(in_buffer[9]*(52))+$signed(in_buffer[10]*(-33))+$signed(in_buffer[11]*(-17))+$signed(in_buffer[12]*(-38))+$signed(in_buffer[13]*(-134))+$signed(in_buffer[14]*(-27))+$signed(in_buffer[15]*(33))+$signed(in_buffer[16]*(38))+$signed(in_buffer[17]*(60))+$signed(in_buffer[18]*(31))+$signed(in_buffer[19]*(-8))+$signed(in_buffer[20]*(-3))+$signed(in_buffer[21]*(23))+$signed(in_buffer[22]*(46))+$signed(in_buffer[23]*(-9))+$signed(in_buffer[24]*(-101));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=$signed(in_buffer[0]*(1))+$signed(in_buffer[1]*(68))+$signed(in_buffer[2]*(48))+$signed(in_buffer[3]*(3))+$signed(in_buffer[4]*(-4))+$signed(in_buffer[5]*(-75))+$signed(in_buffer[6]*(-75))+$signed(in_buffer[7]*(12))+$signed(in_buffer[8]*(48))+$signed(in_buffer[9]*(81))+$signed(in_buffer[10]*(-65))+$signed(in_buffer[11]*(-31))+$signed(in_buffer[12]*(-21))+$signed(in_buffer[13]*(-24))+$signed(in_buffer[14]*(-86))+$signed(in_buffer[15]*(62))+$signed(in_buffer[16]*(27))+$signed(in_buffer[17]*(7))+$signed(in_buffer[18]*(-9))+$signed(in_buffer[19]*(20))+$signed(in_buffer[20]*(65))+$signed(in_buffer[21]*(-24))+$signed(in_buffer[22]*(33))+$signed(in_buffer[23]*(31))+$signed(in_buffer[24]*(67));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=$signed(in_buffer[0]*(-57))+$signed(in_buffer[1]*(-39))+$signed(in_buffer[2]*(-11))+$signed(in_buffer[3]*(4))+$signed(in_buffer[4]*(43))+$signed(in_buffer[5]*(92))+$signed(in_buffer[6]*(67))+$signed(in_buffer[7]*(-8))+$signed(in_buffer[8]*(-67))+$signed(in_buffer[9]*(58))+$signed(in_buffer[10]*(-21))+$signed(in_buffer[11]*(-18))+$signed(in_buffer[12]*(24))+$signed(in_buffer[13]*(25))+$signed(in_buffer[14]*(14))+$signed(in_buffer[15]*(-49))+$signed(in_buffer[16]*(-8))+$signed(in_buffer[17]*(26))+$signed(in_buffer[18]*(-77))+$signed(in_buffer[19]*(-52))+$signed(in_buffer[20]*(-38))+$signed(in_buffer[21]*(11))+$signed(in_buffer[22]*(35))+$signed(in_buffer[23]*(17))+$signed(in_buffer[24]*(33));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=$signed(in_buffer[0]*(64))+$signed(in_buffer[1]*(-120))+$signed(in_buffer[2]*(22))+$signed(in_buffer[3]*(56))+$signed(in_buffer[4]*(16))+$signed(in_buffer[5]*(-91))+$signed(in_buffer[6]*(-4))+$signed(in_buffer[7]*(82))+$signed(in_buffer[8]*(-25))+$signed(in_buffer[9]*(-54))+$signed(in_buffer[10]*(-26))+$signed(in_buffer[11]*(22))+$signed(in_buffer[12]*(18))+$signed(in_buffer[13]*(-25))+$signed(in_buffer[14]*(10))+$signed(in_buffer[15]*(-7))+$signed(in_buffer[16]*(-20))+$signed(in_buffer[17]*(9))+$signed(in_buffer[18]*(28))+$signed(in_buffer[19]*(-178))+$signed(in_buffer[20]*(-6))+$signed(in_buffer[21]*(25))+$signed(in_buffer[22]*(-16))+$signed(in_buffer[23]*(-130))+$signed(in_buffer[24]*(-78));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight10;
assign in_buffer_weight10=$signed(in_buffer[0]*(-33))+$signed(in_buffer[1]*(35))+$signed(in_buffer[2]*(29))+$signed(in_buffer[3]*(-47))+$signed(in_buffer[4]*(-39))+$signed(in_buffer[5]*(-42))+$signed(in_buffer[6]*(-21))+$signed(in_buffer[7]*(-79))+$signed(in_buffer[8]*(33))+$signed(in_buffer[9]*(-29))+$signed(in_buffer[10]*(13))+$signed(in_buffer[11]*(57))+$signed(in_buffer[12]*(52))+$signed(in_buffer[13]*(16))+$signed(in_buffer[14]*(-9))+$signed(in_buffer[15]*(9))+$signed(in_buffer[16]*(17))+$signed(in_buffer[17]*(6))+$signed(in_buffer[18]*(45))+$signed(in_buffer[19]*(-29))+$signed(in_buffer[20]*(0))+$signed(in_buffer[21]*(-22))+$signed(in_buffer[22]*(-5))+$signed(in_buffer[23]*(21))+$signed(in_buffer[24]*(24));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight11;
assign in_buffer_weight11=$signed(in_buffer[0]*(16))+$signed(in_buffer[1]*(85))+$signed(in_buffer[2]*(18))+$signed(in_buffer[3]*(-130))+$signed(in_buffer[4]*(-86))+$signed(in_buffer[5]*(20))+$signed(in_buffer[6]*(-52))+$signed(in_buffer[7]*(3))+$signed(in_buffer[8]*(3))+$signed(in_buffer[9]*(-78))+$signed(in_buffer[10]*(14))+$signed(in_buffer[11]*(-37))+$signed(in_buffer[12]*(59))+$signed(in_buffer[13]*(55))+$signed(in_buffer[14]*(2))+$signed(in_buffer[15]*(45))+$signed(in_buffer[16]*(27))+$signed(in_buffer[17]*(23))+$signed(in_buffer[18]*(-35))+$signed(in_buffer[19]*(-30))+$signed(in_buffer[20]*(-27))+$signed(in_buffer[21]*(-43))+$signed(in_buffer[22]*(-24))+$signed(in_buffer[23]*(-21))+$signed(in_buffer[24]*(-33));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight12;
assign in_buffer_weight12=$signed(in_buffer[0]*(32))+$signed(in_buffer[1]*(2))+$signed(in_buffer[2]*(-62))+$signed(in_buffer[3]*(-9))+$signed(in_buffer[4]*(8))+$signed(in_buffer[5]*(30))+$signed(in_buffer[6]*(97))+$signed(in_buffer[7]*(-34))+$signed(in_buffer[8]*(-5))+$signed(in_buffer[9]*(3))+$signed(in_buffer[10]*(16))+$signed(in_buffer[11]*(54))+$signed(in_buffer[12]*(21))+$signed(in_buffer[13]*(36))+$signed(in_buffer[14]*(-13))+$signed(in_buffer[15]*(-17))+$signed(in_buffer[16]*(0))+$signed(in_buffer[17]*(-36))+$signed(in_buffer[18]*(-40))+$signed(in_buffer[19]*(-28))+$signed(in_buffer[20]*(-64))+$signed(in_buffer[21]*(-11))+$signed(in_buffer[22]*(37))+$signed(in_buffer[23]*(39))+$signed(in_buffer[24]*(23));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight13;
assign in_buffer_weight13=$signed(in_buffer[0]*(-64))+$signed(in_buffer[1]*(-5))+$signed(in_buffer[2]*(53))+$signed(in_buffer[3]*(16))+$signed(in_buffer[4]*(-4))+$signed(in_buffer[5]*(47))+$signed(in_buffer[6]*(36))+$signed(in_buffer[7]*(34))+$signed(in_buffer[8]*(7))+$signed(in_buffer[9]*(43))+$signed(in_buffer[10]*(-7))+$signed(in_buffer[11]*(-17))+$signed(in_buffer[12]*(15))+$signed(in_buffer[13]*(15))+$signed(in_buffer[14]*(-9))+$signed(in_buffer[15]*(3))+$signed(in_buffer[16]*(-1))+$signed(in_buffer[17]*(-67))+$signed(in_buffer[18]*(-16))+$signed(in_buffer[19]*(-47))+$signed(in_buffer[20]*(-14))+$signed(in_buffer[21]*(-5))+$signed(in_buffer[22]*(34))+$signed(in_buffer[23]*(19))+$signed(in_buffer[24]*(11));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight14;
assign in_buffer_weight14=$signed(in_buffer[0]*(4))+$signed(in_buffer[1]*(0))+$signed(in_buffer[2]*(31))+$signed(in_buffer[3]*(23))+$signed(in_buffer[4]*(-28))+$signed(in_buffer[5]*(20))+$signed(in_buffer[6]*(40))+$signed(in_buffer[7]*(-25))+$signed(in_buffer[8]*(27))+$signed(in_buffer[9]*(19))+$signed(in_buffer[10]*(22))+$signed(in_buffer[11]*(-47))+$signed(in_buffer[12]*(-86))+$signed(in_buffer[13]*(87))+$signed(in_buffer[14]*(-45))+$signed(in_buffer[15]*(-15))+$signed(in_buffer[16]*(-37))+$signed(in_buffer[17]*(7))+$signed(in_buffer[18]*(25))+$signed(in_buffer[19]*(-91))+$signed(in_buffer[20]*(23))+$signed(in_buffer[21]*(-28))+$signed(in_buffer[22]*(6))+$signed(in_buffer[23]*(29))+$signed(in_buffer[24]*(87));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight15;
assign in_buffer_weight15=$signed(in_buffer[0]*(-20))+$signed(in_buffer[1]*(16))+$signed(in_buffer[2]*(4))+$signed(in_buffer[3]*(-47))+$signed(in_buffer[4]*(-18))+$signed(in_buffer[5]*(-30))+$signed(in_buffer[6]*(20))+$signed(in_buffer[7]*(9))+$signed(in_buffer[8]*(13))+$signed(in_buffer[9]*(106))+$signed(in_buffer[10]*(14))+$signed(in_buffer[11]*(0))+$signed(in_buffer[12]*(27))+$signed(in_buffer[13]*(-52))+$signed(in_buffer[14]*(-1))+$signed(in_buffer[15]*(-36))+$signed(in_buffer[16]*(-14))+$signed(in_buffer[17]*(56))+$signed(in_buffer[18]*(-94))+$signed(in_buffer[19]*(-75))+$signed(in_buffer[20]*(-37))+$signed(in_buffer[21]*(92))+$signed(in_buffer[22]*(-21))+$signed(in_buffer[23]*(-170))+$signed(in_buffer[24]*(-32));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight16;
assign in_buffer_weight16=$signed(in_buffer[0]*(-11))+$signed(in_buffer[1]*(21))+$signed(in_buffer[2]*(47))+$signed(in_buffer[3]*(14))+$signed(in_buffer[4]*(-30))+$signed(in_buffer[5]*(-21))+$signed(in_buffer[6]*(0))+$signed(in_buffer[7]*(-26))+$signed(in_buffer[8]*(10))+$signed(in_buffer[9]*(10))+$signed(in_buffer[10]*(-19))+$signed(in_buffer[11]*(42))+$signed(in_buffer[12]*(30))+$signed(in_buffer[13]*(-60))+$signed(in_buffer[14]*(45))+$signed(in_buffer[15]*(3))+$signed(in_buffer[16]*(45))+$signed(in_buffer[17]*(-21))+$signed(in_buffer[18]*(40))+$signed(in_buffer[19]*(34))+$signed(in_buffer[20]*(-25))+$signed(in_buffer[21]*(-5))+$signed(in_buffer[22]*(-3))+$signed(in_buffer[23]*(3))+$signed(in_buffer[24]*(-33));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight17;
assign in_buffer_weight17=$signed(in_buffer[0]*(17))+$signed(in_buffer[1]*(-6))+$signed(in_buffer[2]*(10))+$signed(in_buffer[3]*(-4))+$signed(in_buffer[4]*(-4))+$signed(in_buffer[5]*(13))+$signed(in_buffer[6]*(-51))+$signed(in_buffer[7]*(17))+$signed(in_buffer[8]*(-24))+$signed(in_buffer[9]*(23))+$signed(in_buffer[10]*(-22))+$signed(in_buffer[11]*(-1))+$signed(in_buffer[12]*(45))+$signed(in_buffer[13]*(-64))+$signed(in_buffer[14]*(-49))+$signed(in_buffer[15]*(29))+$signed(in_buffer[16]*(-8))+$signed(in_buffer[17]*(18))+$signed(in_buffer[18]*(44))+$signed(in_buffer[19]*(65))+$signed(in_buffer[20]*(6))+$signed(in_buffer[21]*(30))+$signed(in_buffer[22]*(2))+$signed(in_buffer[23]*(33))+$signed(in_buffer[24]*(-31));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight18;
assign in_buffer_weight18=$signed(in_buffer[0]*(26))+$signed(in_buffer[1]*(-45))+$signed(in_buffer[2]*(-6))+$signed(in_buffer[3]*(54))+$signed(in_buffer[4]*(41))+$signed(in_buffer[5]*(-77))+$signed(in_buffer[6]*(-2))+$signed(in_buffer[7]*(-1))+$signed(in_buffer[8]*(-75))+$signed(in_buffer[9]*(-91))+$signed(in_buffer[10]*(53))+$signed(in_buffer[11]*(6))+$signed(in_buffer[12]*(8))+$signed(in_buffer[13]*(43))+$signed(in_buffer[14]*(-15))+$signed(in_buffer[15]*(32))+$signed(in_buffer[16]*(-9))+$signed(in_buffer[17]*(15))+$signed(in_buffer[18]*(71))+$signed(in_buffer[19]*(-20))+$signed(in_buffer[20]*(-31))+$signed(in_buffer[21]*(-3))+$signed(in_buffer[22]*(-28))+$signed(in_buffer[23]*(-67))+$signed(in_buffer[24]*(-6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight19;
assign in_buffer_weight19=$signed(in_buffer[0]*(0))+$signed(in_buffer[1]*(-22))+$signed(in_buffer[2]*(-8))+$signed(in_buffer[3]*(20))+$signed(in_buffer[4]*(-18))+$signed(in_buffer[5]*(-3))+$signed(in_buffer[6]*(21))+$signed(in_buffer[7]*(-1))+$signed(in_buffer[8]*(-6))+$signed(in_buffer[9]*(15))+$signed(in_buffer[10]*(-16))+$signed(in_buffer[11]*(13))+$signed(in_buffer[12]*(-26))+$signed(in_buffer[13]*(-16))+$signed(in_buffer[14]*(18))+$signed(in_buffer[15]*(-14))+$signed(in_buffer[16]*(-22))+$signed(in_buffer[17]*(8))+$signed(in_buffer[18]*(0))+$signed(in_buffer[19]*(-25))+$signed(in_buffer[20]*(10))+$signed(in_buffer[21]*(-24))+$signed(in_buffer[22]*(12))+$signed(in_buffer[23]*(-25))+$signed(in_buffer[24]*(-26));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight20;
assign in_buffer_weight20=$signed(in_buffer[0]*(-15))+$signed(in_buffer[1]*(18))+$signed(in_buffer[2]*(-6))+$signed(in_buffer[3]*(8))+$signed(in_buffer[4]*(-5))+$signed(in_buffer[5]*(0))+$signed(in_buffer[6]*(-11))+$signed(in_buffer[7]*(19))+$signed(in_buffer[8]*(-2))+$signed(in_buffer[9]*(7))+$signed(in_buffer[10]*(-27))+$signed(in_buffer[11]*(1))+$signed(in_buffer[12]*(-1))+$signed(in_buffer[13]*(-27))+$signed(in_buffer[14]*(-10))+$signed(in_buffer[15]*(-6))+$signed(in_buffer[16]*(-5))+$signed(in_buffer[17]*(-21))+$signed(in_buffer[18]*(3))+$signed(in_buffer[19]*(17))+$signed(in_buffer[20]*(-17))+$signed(in_buffer[21]*(-9))+$signed(in_buffer[22]*(13))+$signed(in_buffer[23]*(-10))+$signed(in_buffer[24]*(-5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight21;
assign in_buffer_weight21=$signed(in_buffer[0]*(-56))+$signed(in_buffer[1]*(22))+$signed(in_buffer[2]*(10))+$signed(in_buffer[3]*(3))+$signed(in_buffer[4]*(19))+$signed(in_buffer[5]*(43))+$signed(in_buffer[6]*(-4))+$signed(in_buffer[7]*(-28))+$signed(in_buffer[8]*(-21))+$signed(in_buffer[9]*(36))+$signed(in_buffer[10]*(-2))+$signed(in_buffer[11]*(73))+$signed(in_buffer[12]*(65))+$signed(in_buffer[13]*(-33))+$signed(in_buffer[14]*(-71))+$signed(in_buffer[15]*(-119))+$signed(in_buffer[16]*(-90))+$signed(in_buffer[17]*(-43))+$signed(in_buffer[18]*(48))+$signed(in_buffer[19]*(17))+$signed(in_buffer[20]*(73))+$signed(in_buffer[21]*(59))+$signed(in_buffer[22]*(-1))+$signed(in_buffer[23]*(6))+$signed(in_buffer[24]*(58));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight22;
assign in_buffer_weight22=$signed(in_buffer[0]*(17))+$signed(in_buffer[1]*(65))+$signed(in_buffer[2]*(112))+$signed(in_buffer[3]*(51))+$signed(in_buffer[4]*(-11))+$signed(in_buffer[5]*(-8))+$signed(in_buffer[6]*(-44))+$signed(in_buffer[7]*(-33))+$signed(in_buffer[8]*(22))+$signed(in_buffer[9]*(17))+$signed(in_buffer[10]*(-5))+$signed(in_buffer[11]*(-40))+$signed(in_buffer[12]*(-34))+$signed(in_buffer[13]*(64))+$signed(in_buffer[14]*(-110))+$signed(in_buffer[15]*(10))+$signed(in_buffer[16]*(-27))+$signed(in_buffer[17]*(-23))+$signed(in_buffer[18]*(2))+$signed(in_buffer[19]*(-112))+$signed(in_buffer[20]*(50))+$signed(in_buffer[21]*(31))+$signed(in_buffer[22]*(45))+$signed(in_buffer[23]*(-9))+$signed(in_buffer[24]*(10));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight23;
assign in_buffer_weight23=$signed(in_buffer[0]*(85))+$signed(in_buffer[1]*(-45))+$signed(in_buffer[2]*(-8))+$signed(in_buffer[3]*(35))+$signed(in_buffer[4]*(-60))+$signed(in_buffer[5]*(-60))+$signed(in_buffer[6]*(-105))+$signed(in_buffer[7]*(17))+$signed(in_buffer[8]*(12))+$signed(in_buffer[9]*(-76))+$signed(in_buffer[10]*(-4))+$signed(in_buffer[11]*(44))+$signed(in_buffer[12]*(28))+$signed(in_buffer[13]*(-14))+$signed(in_buffer[14]*(33))+$signed(in_buffer[15]*(78))+$signed(in_buffer[16]*(-45))+$signed(in_buffer[17]*(29))+$signed(in_buffer[18]*(39))+$signed(in_buffer[19]*(51))+$signed(in_buffer[20]*(-8))+$signed(in_buffer[21]*(-13))+$signed(in_buffer[22]*(-31))+$signed(in_buffer[23]*(46))+$signed(in_buffer[24]*(-57));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight24;
assign in_buffer_weight24=$signed(in_buffer[0]*(10))+$signed(in_buffer[1]*(41))+$signed(in_buffer[2]*(51))+$signed(in_buffer[3]*(30))+$signed(in_buffer[4]*(-33))+$signed(in_buffer[5]*(-41))+$signed(in_buffer[6]*(-40))+$signed(in_buffer[7]*(-20))+$signed(in_buffer[8]*(2))+$signed(in_buffer[9]*(36))+$signed(in_buffer[10]*(18))+$signed(in_buffer[11]*(51))+$signed(in_buffer[12]*(-5))+$signed(in_buffer[13]*(-8))+$signed(in_buffer[14]*(-2))+$signed(in_buffer[15]*(46))+$signed(in_buffer[16]*(82))+$signed(in_buffer[17]*(-65))+$signed(in_buffer[18]*(-43))+$signed(in_buffer[19]*(13))+$signed(in_buffer[20]*(44))+$signed(in_buffer[21]*(63))+$signed(in_buffer[22]*(-42))+$signed(in_buffer[23]*(-13))+$signed(in_buffer[24]*(-33));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight25;
assign in_buffer_weight25=$signed(in_buffer[0]*(34))+$signed(in_buffer[1]*(37))+$signed(in_buffer[2]*(19))+$signed(in_buffer[3]*(-36))+$signed(in_buffer[4]*(-22))+$signed(in_buffer[5]*(-16))+$signed(in_buffer[6]*(15))+$signed(in_buffer[7]*(-67))+$signed(in_buffer[8]*(16))+$signed(in_buffer[9]*(20))+$signed(in_buffer[10]*(8))+$signed(in_buffer[11]*(19))+$signed(in_buffer[12]*(67))+$signed(in_buffer[13]*(15))+$signed(in_buffer[14]*(5))+$signed(in_buffer[15]*(5))+$signed(in_buffer[16]*(14))+$signed(in_buffer[17]*(-50))+$signed(in_buffer[18]*(4))+$signed(in_buffer[19]*(-54))+$signed(in_buffer[20]*(-30))+$signed(in_buffer[21]*(13))+$signed(in_buffer[22]*(61))+$signed(in_buffer[23]*(18))+$signed(in_buffer[24]*(-60));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight26;
assign in_buffer_weight26=$signed(in_buffer[0]*(19))+$signed(in_buffer[1]*(7))+$signed(in_buffer[2]*(-69))+$signed(in_buffer[3]*(-108))+$signed(in_buffer[4]*(-54))+$signed(in_buffer[5]*(1))+$signed(in_buffer[6]*(-18))+$signed(in_buffer[7]*(58))+$signed(in_buffer[8]*(22))+$signed(in_buffer[9]*(33))+$signed(in_buffer[10]*(-31))+$signed(in_buffer[11]*(-15))+$signed(in_buffer[12]*(29))+$signed(in_buffer[13]*(-30))+$signed(in_buffer[14]*(16))+$signed(in_buffer[15]*(25))+$signed(in_buffer[16]*(41))+$signed(in_buffer[17]*(85))+$signed(in_buffer[18]*(40))+$signed(in_buffer[19]*(-6))+$signed(in_buffer[20]*(-79))+$signed(in_buffer[21]*(-38))+$signed(in_buffer[22]*(-68))+$signed(in_buffer[23]*(-136))+$signed(in_buffer[24]*(-55));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight27;
assign in_buffer_weight27=$signed(in_buffer[0]*(-32))+$signed(in_buffer[1]*(-2))+$signed(in_buffer[2]*(1))+$signed(in_buffer[3]*(99))+$signed(in_buffer[4]*(130))+$signed(in_buffer[5]*(-5))+$signed(in_buffer[6]*(23))+$signed(in_buffer[7]*(14))+$signed(in_buffer[8]*(-81))+$signed(in_buffer[9]*(-118))+$signed(in_buffer[10]*(10))+$signed(in_buffer[11]*(-56))+$signed(in_buffer[12]*(3))+$signed(in_buffer[13]*(-5))+$signed(in_buffer[14]*(-44))+$signed(in_buffer[15]*(25))+$signed(in_buffer[16]*(12))+$signed(in_buffer[17]*(52))+$signed(in_buffer[18]*(-11))+$signed(in_buffer[19]*(22))+$signed(in_buffer[20]*(-40))+$signed(in_buffer[21]*(-45))+$signed(in_buffer[22]*(-6))+$signed(in_buffer[23]*(45))+$signed(in_buffer[24]*(26));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight28;
assign in_buffer_weight28=$signed(in_buffer[0]*(0))+$signed(in_buffer[1]*(24))+$signed(in_buffer[2]*(3))+$signed(in_buffer[3]*(33))+$signed(in_buffer[4]*(39))+$signed(in_buffer[5]*(18))+$signed(in_buffer[6]*(-61))+$signed(in_buffer[7]*(-33))+$signed(in_buffer[8]*(61))+$signed(in_buffer[9]*(-22))+$signed(in_buffer[10]*(0))+$signed(in_buffer[11]*(42))+$signed(in_buffer[12]*(60))+$signed(in_buffer[13]*(75))+$signed(in_buffer[14]*(8))+$signed(in_buffer[15]*(-1))+$signed(in_buffer[16]*(-58))+$signed(in_buffer[17]*(-44))+$signed(in_buffer[18]*(-41))+$signed(in_buffer[19]*(-17))+$signed(in_buffer[20]*(8))+$signed(in_buffer[21]*(-52))+$signed(in_buffer[22]*(-3))+$signed(in_buffer[23]*(2))+$signed(in_buffer[24]*(15));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight29;
assign in_buffer_weight29=$signed(in_buffer[0]*(-27))+$signed(in_buffer[1]*(-10))+$signed(in_buffer[2]*(43))+$signed(in_buffer[3]*(-48))+$signed(in_buffer[4]*(-54))+$signed(in_buffer[5]*(-56))+$signed(in_buffer[6]*(23))+$signed(in_buffer[7]*(5))+$signed(in_buffer[8]*(7))+$signed(in_buffer[9]*(-1))+$signed(in_buffer[10]*(-30))+$signed(in_buffer[11]*(16))+$signed(in_buffer[12]*(-15))+$signed(in_buffer[13]*(36))+$signed(in_buffer[14]*(-16))+$signed(in_buffer[15]*(-102))+$signed(in_buffer[16]*(31))+$signed(in_buffer[17]*(5))+$signed(in_buffer[18]*(12))+$signed(in_buffer[19]*(-38))+$signed(in_buffer[20]*(-298))+$signed(in_buffer[21]*(-106))+$signed(in_buffer[22]*(43))+$signed(in_buffer[23]*(-4))+$signed(in_buffer[24]*(-23));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight30;
assign in_buffer_weight30=$signed(in_buffer[0]*(21))+$signed(in_buffer[1]*(-1))+$signed(in_buffer[2]*(-16))+$signed(in_buffer[3]*(-11))+$signed(in_buffer[4]*(-51))+$signed(in_buffer[5]*(52))+$signed(in_buffer[6]*(39))+$signed(in_buffer[7]*(-62))+$signed(in_buffer[8]*(-29))+$signed(in_buffer[9]*(40))+$signed(in_buffer[10]*(-3))+$signed(in_buffer[11]*(-98))+$signed(in_buffer[12]*(36))+$signed(in_buffer[13]*(3))+$signed(in_buffer[14]*(39))+$signed(in_buffer[15]*(-60))+$signed(in_buffer[16]*(20))+$signed(in_buffer[17]*(108))+$signed(in_buffer[18]*(-8))+$signed(in_buffer[19]*(20))+$signed(in_buffer[20]*(8))+$signed(in_buffer[21]*(-28))+$signed(in_buffer[22]*(15))+$signed(in_buffer[23]*(6))+$signed(in_buffer[24]*(11));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight31;
assign in_buffer_weight31=$signed(in_buffer[0]*(8))+$signed(in_buffer[1]*(-26))+$signed(in_buffer[2]*(-10))+$signed(in_buffer[3]*(31))+$signed(in_buffer[4]*(83))+$signed(in_buffer[5]*(65))+$signed(in_buffer[6]*(25))+$signed(in_buffer[7]*(68))+$signed(in_buffer[8]*(-16))+$signed(in_buffer[9]*(4))+$signed(in_buffer[10]*(-30))+$signed(in_buffer[11]*(-53))+$signed(in_buffer[12]*(-55))+$signed(in_buffer[13]*(-44))+$signed(in_buffer[14]*(-27))+$signed(in_buffer[15]*(1))+$signed(in_buffer[16]*(9))+$signed(in_buffer[17]*(26))+$signed(in_buffer[18]*(10))+$signed(in_buffer[19]*(31))+$signed(in_buffer[20]*(21))+$signed(in_buffer[21]*(14))+$signed(in_buffer[22]*(19))+$signed(in_buffer[23]*(45))+$signed(in_buffer[24]*(-62));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight32;
assign in_buffer_weight32=$signed(in_buffer[0]*(10))+$signed(in_buffer[1]*(-23))+$signed(in_buffer[2]*(-12))+$signed(in_buffer[3]*(4))+$signed(in_buffer[4]*(-23))+$signed(in_buffer[5]*(-11))+$signed(in_buffer[6]*(-14))+$signed(in_buffer[7]*(-1))+$signed(in_buffer[8]*(0))+$signed(in_buffer[9]*(-14))+$signed(in_buffer[10]*(-4))+$signed(in_buffer[11]*(-5))+$signed(in_buffer[12]*(-5))+$signed(in_buffer[13]*(-11))+$signed(in_buffer[14]*(24))+$signed(in_buffer[15]*(20))+$signed(in_buffer[16]*(-12))+$signed(in_buffer[17]*(-20))+$signed(in_buffer[18]*(-4))+$signed(in_buffer[19]*(1))+$signed(in_buffer[20]*(7))+$signed(in_buffer[21]*(-13))+$signed(in_buffer[22]*(9))+$signed(in_buffer[23]*(-10))+$signed(in_buffer[24]*(25));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight33;
assign in_buffer_weight33=$signed(in_buffer[0]*(-6))+$signed(in_buffer[1]*(-16))+$signed(in_buffer[2]*(12))+$signed(in_buffer[3]*(26))+$signed(in_buffer[4]*(-116))+$signed(in_buffer[5]*(11))+$signed(in_buffer[6]*(-59))+$signed(in_buffer[7]*(47))+$signed(in_buffer[8]*(21))+$signed(in_buffer[9]*(-228))+$signed(in_buffer[10]*(59))+$signed(in_buffer[11]*(-5))+$signed(in_buffer[12]*(27))+$signed(in_buffer[13]*(-11))+$signed(in_buffer[14]*(54))+$signed(in_buffer[15]*(-27))+$signed(in_buffer[16]*(-4))+$signed(in_buffer[17]*(69))+$signed(in_buffer[18]*(-83))+$signed(in_buffer[19]*(33))+$signed(in_buffer[20]*(-84))+$signed(in_buffer[21]*(-21))+$signed(in_buffer[22]*(10))+$signed(in_buffer[23]*(-2))+$signed(in_buffer[24]*(-79));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight34;
assign in_buffer_weight34=$signed(in_buffer[0]*(-22))+$signed(in_buffer[1]*(-17))+$signed(in_buffer[2]*(27))+$signed(in_buffer[3]*(17))+$signed(in_buffer[4]*(-6))+$signed(in_buffer[5]*(-16))+$signed(in_buffer[6]*(29))+$signed(in_buffer[7]*(-26))+$signed(in_buffer[8]*(-20))+$signed(in_buffer[9]*(36))+$signed(in_buffer[10]*(49))+$signed(in_buffer[11]*(28))+$signed(in_buffer[12]*(-1))+$signed(in_buffer[13]*(-69))+$signed(in_buffer[14]*(56))+$signed(in_buffer[15]*(10))+$signed(in_buffer[16]*(46))+$signed(in_buffer[17]*(-11))+$signed(in_buffer[18]*(53))+$signed(in_buffer[19]*(26))+$signed(in_buffer[20]*(-37))+$signed(in_buffer[21]*(39))+$signed(in_buffer[22]*(-2))+$signed(in_buffer[23]*(-37))+$signed(in_buffer[24]*(-112));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight35;
assign in_buffer_weight35=$signed(in_buffer[0]*(-30))+$signed(in_buffer[1]*(-8))+$signed(in_buffer[2]*(-6))+$signed(in_buffer[3]*(-57))+$signed(in_buffer[4]*(-11))+$signed(in_buffer[5]*(-6))+$signed(in_buffer[6]*(29))+$signed(in_buffer[7]*(68))+$signed(in_buffer[8]*(37))+$signed(in_buffer[9]*(-163))+$signed(in_buffer[10]*(-2))+$signed(in_buffer[11]*(-19))+$signed(in_buffer[12]*(14))+$signed(in_buffer[13]*(-64))+$signed(in_buffer[14]*(-214))+$signed(in_buffer[15]*(-6))+$signed(in_buffer[16]*(19))+$signed(in_buffer[17]*(24))+$signed(in_buffer[18]*(-52))+$signed(in_buffer[19]*(141))+$signed(in_buffer[20]*(16))+$signed(in_buffer[21]*(-6))+$signed(in_buffer[22]*(-12))+$signed(in_buffer[23]*(52))+$signed(in_buffer[24]*(-37));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight36;
assign in_buffer_weight36=$signed(in_buffer[0]*(-55))+$signed(in_buffer[1]*(29))+$signed(in_buffer[2]*(5))+$signed(in_buffer[3]*(1))+$signed(in_buffer[4]*(49))+$signed(in_buffer[5]*(-29))+$signed(in_buffer[6]*(23))+$signed(in_buffer[7]*(-23))+$signed(in_buffer[8]*(0))+$signed(in_buffer[9]*(-22))+$signed(in_buffer[10]*(53))+$signed(in_buffer[11]*(25))+$signed(in_buffer[12]*(48))+$signed(in_buffer[13]*(69))+$signed(in_buffer[14]*(-1))+$signed(in_buffer[15]*(-128))+$signed(in_buffer[16]*(-75))+$signed(in_buffer[17]*(0))+$signed(in_buffer[18]*(-51))+$signed(in_buffer[19]*(-9))+$signed(in_buffer[20]*(-10))+$signed(in_buffer[21]*(79))+$signed(in_buffer[22]*(-47))+$signed(in_buffer[23]*(-238))+$signed(in_buffer[24]*(52));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight37;
assign in_buffer_weight37=$signed(in_buffer[0]*(3))+$signed(in_buffer[1]*(-11))+$signed(in_buffer[2]*(37))+$signed(in_buffer[3]*(9))+$signed(in_buffer[4]*(-82))+$signed(in_buffer[5]*(1))+$signed(in_buffer[6]*(-26))+$signed(in_buffer[7]*(28))+$signed(in_buffer[8]*(24))+$signed(in_buffer[9]*(35))+$signed(in_buffer[10]*(16))+$signed(in_buffer[11]*(-44))+$signed(in_buffer[12]*(27))+$signed(in_buffer[13]*(-27))+$signed(in_buffer[14]*(21))+$signed(in_buffer[15]*(-5))+$signed(in_buffer[16]*(17))+$signed(in_buffer[17]*(-41))+$signed(in_buffer[18]*(53))+$signed(in_buffer[19]*(20))+$signed(in_buffer[20]*(-7))+$signed(in_buffer[21]*(58))+$signed(in_buffer[22]*(51))+$signed(in_buffer[23]*(7))+$signed(in_buffer[24]*(-63));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight38;
assign in_buffer_weight38=$signed(in_buffer[0]*(-23))+$signed(in_buffer[1]*(-29))+$signed(in_buffer[2]*(38))+$signed(in_buffer[3]*(-2))+$signed(in_buffer[4]*(-49))+$signed(in_buffer[5]*(53))+$signed(in_buffer[6]*(20))+$signed(in_buffer[7]*(-16))+$signed(in_buffer[8]*(21))+$signed(in_buffer[9]*(40))+$signed(in_buffer[10]*(-27))+$signed(in_buffer[11]*(-18))+$signed(in_buffer[12]*(9))+$signed(in_buffer[13]*(11))+$signed(in_buffer[14]*(-10))+$signed(in_buffer[15]*(-55))+$signed(in_buffer[16]*(50))+$signed(in_buffer[17]*(-48))+$signed(in_buffer[18]*(-9))+$signed(in_buffer[19]*(-12))+$signed(in_buffer[20]*(-28))+$signed(in_buffer[21]*(29))+$signed(in_buffer[22]*(58))+$signed(in_buffer[23]*(3))+$signed(in_buffer[24]*(21));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight39;
assign in_buffer_weight39=$signed(in_buffer[0]*(-256))+$signed(in_buffer[1]*(69))+$signed(in_buffer[2]*(21))+$signed(in_buffer[3]*(-98))+$signed(in_buffer[4]*(54))+$signed(in_buffer[5]*(-117))+$signed(in_buffer[6]*(67))+$signed(in_buffer[7]*(-54))+$signed(in_buffer[8]*(-31))+$signed(in_buffer[9]*(29))+$signed(in_buffer[10]*(-35))+$signed(in_buffer[11]*(25))+$signed(in_buffer[12]*(-17))+$signed(in_buffer[13]*(7))+$signed(in_buffer[14]*(11))+$signed(in_buffer[15]*(13))+$signed(in_buffer[16]*(30))+$signed(in_buffer[17]*(11))+$signed(in_buffer[18]*(19))+$signed(in_buffer[19]*(24))+$signed(in_buffer[20]*(-32))+$signed(in_buffer[21]*(31))+$signed(in_buffer[22]*(8))+$signed(in_buffer[23]*(17))+$signed(in_buffer[24]*(-53));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight40;
assign in_buffer_weight40=$signed(in_buffer[0]*(-11))+$signed(in_buffer[1]*(-15))+$signed(in_buffer[2]*(22))+$signed(in_buffer[3]*(8))+$signed(in_buffer[4]*(-22))+$signed(in_buffer[5]*(22))+$signed(in_buffer[6]*(-9))+$signed(in_buffer[7]*(-22))+$signed(in_buffer[8]*(-16))+$signed(in_buffer[9]*(-15))+$signed(in_buffer[10]*(-10))+$signed(in_buffer[11]*(11))+$signed(in_buffer[12]*(-15))+$signed(in_buffer[13]*(-14))+$signed(in_buffer[14]*(-17))+$signed(in_buffer[15]*(-9))+$signed(in_buffer[16]*(13))+$signed(in_buffer[17]*(5))+$signed(in_buffer[18]*(-21))+$signed(in_buffer[19]*(24))+$signed(in_buffer[20]*(7))+$signed(in_buffer[21]*(9))+$signed(in_buffer[22]*(-9))+$signed(in_buffer[23]*(14))+$signed(in_buffer[24]*(-17));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight41;
assign in_buffer_weight41=$signed(in_buffer[0]*(44))+$signed(in_buffer[1]*(-33))+$signed(in_buffer[2]*(-20))+$signed(in_buffer[3]*(13))+$signed(in_buffer[4]*(24))+$signed(in_buffer[5]*(-8))+$signed(in_buffer[6]*(41))+$signed(in_buffer[7]*(25))+$signed(in_buffer[8]*(-7))+$signed(in_buffer[9]*(-27))+$signed(in_buffer[10]*(53))+$signed(in_buffer[11]*(18))+$signed(in_buffer[12]*(-81))+$signed(in_buffer[13]*(40))+$signed(in_buffer[14]*(-14))+$signed(in_buffer[15]*(14))+$signed(in_buffer[16]*(-30))+$signed(in_buffer[17]*(35))+$signed(in_buffer[18]*(53))+$signed(in_buffer[19]*(-32))+$signed(in_buffer[20]*(-22))+$signed(in_buffer[21]*(-31))+$signed(in_buffer[22]*(49))+$signed(in_buffer[23]*(9))+$signed(in_buffer[24]*(-20));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight42;
assign in_buffer_weight42=$signed(in_buffer[0]*(39))+$signed(in_buffer[1]*(-32))+$signed(in_buffer[2]*(23))+$signed(in_buffer[3]*(-58))+$signed(in_buffer[4]*(-129))+$signed(in_buffer[5]*(-27))+$signed(in_buffer[6]*(-14))+$signed(in_buffer[7]*(112))+$signed(in_buffer[8]*(-71))+$signed(in_buffer[9]*(-115))+$signed(in_buffer[10]*(3))+$signed(in_buffer[11]*(43))+$signed(in_buffer[12]*(13))+$signed(in_buffer[13]*(-20))+$signed(in_buffer[14]*(97))+$signed(in_buffer[15]*(31))+$signed(in_buffer[16]*(-40))+$signed(in_buffer[17]*(0))+$signed(in_buffer[18]*(-9))+$signed(in_buffer[19]*(-7))+$signed(in_buffer[20]*(-5))+$signed(in_buffer[21]*(-30))+$signed(in_buffer[22]*(49))+$signed(in_buffer[23]*(-10))+$signed(in_buffer[24]*(-68));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight43;
assign in_buffer_weight43=$signed(in_buffer[0]*(-74))+$signed(in_buffer[1]*(-13))+$signed(in_buffer[2]*(64))+$signed(in_buffer[3]*(54))+$signed(in_buffer[4]*(-72))+$signed(in_buffer[5]*(28))+$signed(in_buffer[6]*(-45))+$signed(in_buffer[7]*(-77))+$signed(in_buffer[8]*(69))+$signed(in_buffer[9]*(60))+$signed(in_buffer[10]*(27))+$signed(in_buffer[11]*(22))+$signed(in_buffer[12]*(-31))+$signed(in_buffer[13]*(23))+$signed(in_buffer[14]*(-36))+$signed(in_buffer[15]*(-7))+$signed(in_buffer[16]*(14))+$signed(in_buffer[17]*(13))+$signed(in_buffer[18]*(11))+$signed(in_buffer[19]*(-71))+$signed(in_buffer[20]*(0))+$signed(in_buffer[21]*(-3))+$signed(in_buffer[22]*(9))+$signed(in_buffer[23]*(9))+$signed(in_buffer[24]*(71));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight44;
assign in_buffer_weight44=$signed(in_buffer[0]*(0))+$signed(in_buffer[1]*(0))+$signed(in_buffer[2]*(-16))+$signed(in_buffer[3]*(16))+$signed(in_buffer[4]*(6))+$signed(in_buffer[5]*(77))+$signed(in_buffer[6]*(8))+$signed(in_buffer[7]*(25))+$signed(in_buffer[8]*(35))+$signed(in_buffer[9]*(-40))+$signed(in_buffer[10]*(-85))+$signed(in_buffer[11]*(-103))+$signed(in_buffer[12]*(76))+$signed(in_buffer[13]*(0))+$signed(in_buffer[14]*(-33))+$signed(in_buffer[15]*(-48))+$signed(in_buffer[16]*(-20))+$signed(in_buffer[17]*(13))+$signed(in_buffer[18]*(-8))+$signed(in_buffer[19]*(40))+$signed(in_buffer[20]*(87))+$signed(in_buffer[21]*(28))+$signed(in_buffer[22]*(-5))+$signed(in_buffer[23]*(32))+$signed(in_buffer[24]*(29));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight45;
assign in_buffer_weight45=$signed(in_buffer[0]*(-67))+$signed(in_buffer[1]*(-3))+$signed(in_buffer[2]*(13))+$signed(in_buffer[3]*(27))+$signed(in_buffer[4]*(24))+$signed(in_buffer[5]*(21))+$signed(in_buffer[6]*(69))+$signed(in_buffer[7]*(-15))+$signed(in_buffer[8]*(-57))+$signed(in_buffer[9]*(6))+$signed(in_buffer[10]*(-55))+$signed(in_buffer[11]*(14))+$signed(in_buffer[12]*(14))+$signed(in_buffer[13]*(-77))+$signed(in_buffer[14]*(20))+$signed(in_buffer[15]*(15))+$signed(in_buffer[16]*(20))+$signed(in_buffer[17]*(-53))+$signed(in_buffer[18]*(39))+$signed(in_buffer[19]*(-12))+$signed(in_buffer[20]*(14))+$signed(in_buffer[21]*(27))+$signed(in_buffer[22]*(45))+$signed(in_buffer[23]*(23))+$signed(in_buffer[24]*(-94));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight46;
assign in_buffer_weight46=$signed(in_buffer[0]*(-217))+$signed(in_buffer[1]*(-96))+$signed(in_buffer[2]*(43))+$signed(in_buffer[3]*(41))+$signed(in_buffer[4]*(-23))+$signed(in_buffer[5]*(-43))+$signed(in_buffer[6]*(3))+$signed(in_buffer[7]*(-34))+$signed(in_buffer[8]*(-22))+$signed(in_buffer[9]*(-1))+$signed(in_buffer[10]*(2))+$signed(in_buffer[11]*(29))+$signed(in_buffer[12]*(56))+$signed(in_buffer[13]*(54))+$signed(in_buffer[14]*(-5))+$signed(in_buffer[15]*(-24))+$signed(in_buffer[16]*(16))+$signed(in_buffer[17]*(-44))+$signed(in_buffer[18]*(-46))+$signed(in_buffer[19]*(23))+$signed(in_buffer[20]*(-52))+$signed(in_buffer[21]*(43))+$signed(in_buffer[22]*(-12))+$signed(in_buffer[23]*(-19))+$signed(in_buffer[24]*(18));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight47;
assign in_buffer_weight47=$signed(in_buffer[0]*(147))+$signed(in_buffer[1]*(83))+$signed(in_buffer[2]*(-37))+$signed(in_buffer[3]*(-16))+$signed(in_buffer[4]*(-22))+$signed(in_buffer[5]*(-31))+$signed(in_buffer[6]*(34))+$signed(in_buffer[7]*(-22))+$signed(in_buffer[8]*(1))+$signed(in_buffer[9]*(-28))+$signed(in_buffer[10]*(44))+$signed(in_buffer[11]*(28))+$signed(in_buffer[12]*(-29))+$signed(in_buffer[13]*(60))+$signed(in_buffer[14]*(53))+$signed(in_buffer[15]*(-71))+$signed(in_buffer[16]*(29))+$signed(in_buffer[17]*(25))+$signed(in_buffer[18]*(0))+$signed(in_buffer[19]*(-22))+$signed(in_buffer[20]*(-87))+$signed(in_buffer[21]*(-23))+$signed(in_buffer[22]*(14))+$signed(in_buffer[23]*(-15))+$signed(in_buffer[24]*(27));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight48;
assign in_buffer_weight48=$signed(in_buffer[0]*(-11))+$signed(in_buffer[1]*(4))+$signed(in_buffer[2]*(-25))+$signed(in_buffer[3]*(-27))+$signed(in_buffer[4]*(5))+$signed(in_buffer[5]*(-26))+$signed(in_buffer[6]*(-20))+$signed(in_buffer[7]*(14))+$signed(in_buffer[8]*(-1))+$signed(in_buffer[9]*(-8))+$signed(in_buffer[10]*(-24))+$signed(in_buffer[11]*(-20))+$signed(in_buffer[12]*(16))+$signed(in_buffer[13]*(0))+$signed(in_buffer[14]*(-2))+$signed(in_buffer[15]*(-4))+$signed(in_buffer[16]*(-29))+$signed(in_buffer[17]*(-19))+$signed(in_buffer[18]*(10))+$signed(in_buffer[19]*(-29))+$signed(in_buffer[20]*(10))+$signed(in_buffer[21]*(11))+$signed(in_buffer[22]*(-15))+$signed(in_buffer[23]*(-3))+$signed(in_buffer[24]*(10));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight49;
assign in_buffer_weight49=$signed(in_buffer[0]*(8))+$signed(in_buffer[1]*(12))+$signed(in_buffer[2]*(-40))+$signed(in_buffer[3]*(7))+$signed(in_buffer[4]*(35))+$signed(in_buffer[5]*(8))+$signed(in_buffer[6]*(4))+$signed(in_buffer[7]*(-11))+$signed(in_buffer[8]*(49))+$signed(in_buffer[9]*(11))+$signed(in_buffer[10]*(-62))+$signed(in_buffer[11]*(-5))+$signed(in_buffer[12]*(-51))+$signed(in_buffer[13]*(8))+$signed(in_buffer[14]*(-105))+$signed(in_buffer[15]*(-53))+$signed(in_buffer[16]*(77))+$signed(in_buffer[17]*(1))+$signed(in_buffer[18]*(-15))+$signed(in_buffer[19]*(13))+$signed(in_buffer[20]*(-109))+$signed(in_buffer[21]*(33))+$signed(in_buffer[22]*(41))+$signed(in_buffer[23]*(43))+$signed(in_buffer[24]*(41));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight50;
assign in_buffer_weight50=$signed(in_buffer[0]*(-62))+$signed(in_buffer[1]*(-6))+$signed(in_buffer[2]*(28))+$signed(in_buffer[3]*(-54))+$signed(in_buffer[4]*(-75))+$signed(in_buffer[5]*(-10))+$signed(in_buffer[6]*(-2))+$signed(in_buffer[7]*(43))+$signed(in_buffer[8]*(37))+$signed(in_buffer[9]*(-10))+$signed(in_buffer[10]*(50))+$signed(in_buffer[11]*(-30))+$signed(in_buffer[12]*(-3))+$signed(in_buffer[13]*(38))+$signed(in_buffer[14]*(-10))+$signed(in_buffer[15]*(61))+$signed(in_buffer[16]*(-16))+$signed(in_buffer[17]*(-67))+$signed(in_buffer[18]*(-6))+$signed(in_buffer[19]*(-43))+$signed(in_buffer[20]*(50))+$signed(in_buffer[21]*(30))+$signed(in_buffer[22]*(8))+$signed(in_buffer[23]*(0))+$signed(in_buffer[24]*(-46));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight51;
assign in_buffer_weight51=$signed(in_buffer[0]*(21))+$signed(in_buffer[1]*(49))+$signed(in_buffer[2]*(56))+$signed(in_buffer[3]*(48))+$signed(in_buffer[4]*(48))+$signed(in_buffer[5]*(47))+$signed(in_buffer[6]*(-69))+$signed(in_buffer[7]*(-15))+$signed(in_buffer[8]*(9))+$signed(in_buffer[9]*(-109))+$signed(in_buffer[10]*(-15))+$signed(in_buffer[11]*(-55))+$signed(in_buffer[12]*(22))+$signed(in_buffer[13]*(9))+$signed(in_buffer[14]*(50))+$signed(in_buffer[15]*(-48))+$signed(in_buffer[16]*(25))+$signed(in_buffer[17]*(23))+$signed(in_buffer[18]*(-14))+$signed(in_buffer[19]*(33))+$signed(in_buffer[20]*(7))+$signed(in_buffer[21]*(-16))+$signed(in_buffer[22]*(5))+$signed(in_buffer[23]*(-61))+$signed(in_buffer[24]*(-59));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight52;
assign in_buffer_weight52=$signed(in_buffer[0]*(-171))+$signed(in_buffer[1]*(-12))+$signed(in_buffer[2]*(74))+$signed(in_buffer[3]*(-11))+$signed(in_buffer[4]*(-121))+$signed(in_buffer[5]*(-69))+$signed(in_buffer[6]*(1))+$signed(in_buffer[7]*(7))+$signed(in_buffer[8]*(-35))+$signed(in_buffer[9]*(3))+$signed(in_buffer[10]*(17))+$signed(in_buffer[11]*(72))+$signed(in_buffer[12]*(-62))+$signed(in_buffer[13]*(-1))+$signed(in_buffer[14]*(4))+$signed(in_buffer[15]*(-7))+$signed(in_buffer[16]*(20))+$signed(in_buffer[17]*(7))+$signed(in_buffer[18]*(22))+$signed(in_buffer[19]*(37))+$signed(in_buffer[20]*(-9))+$signed(in_buffer[21]*(53))+$signed(in_buffer[22]*(-34))+$signed(in_buffer[23]*(4))+$signed(in_buffer[24]*(-19));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight53;
assign in_buffer_weight53=$signed(in_buffer[0]*(-3))+$signed(in_buffer[1]*(14))+$signed(in_buffer[2]*(-38))+$signed(in_buffer[3]*(-2))+$signed(in_buffer[4]*(80))+$signed(in_buffer[5]*(-58))+$signed(in_buffer[6]*(2))+$signed(in_buffer[7]*(47))+$signed(in_buffer[8]*(54))+$signed(in_buffer[9]*(-38))+$signed(in_buffer[10]*(1))+$signed(in_buffer[11]*(0))+$signed(in_buffer[12]*(40))+$signed(in_buffer[13]*(-5))+$signed(in_buffer[14]*(-21))+$signed(in_buffer[15]*(3))+$signed(in_buffer[16]*(-52))+$signed(in_buffer[17]*(0))+$signed(in_buffer[18]*(22))+$signed(in_buffer[19]*(-45))+$signed(in_buffer[20]*(10))+$signed(in_buffer[21]*(2))+$signed(in_buffer[22]*(47))+$signed(in_buffer[23]*(0))+$signed(in_buffer[24]*(-280));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight54;
assign in_buffer_weight54=$signed(in_buffer[0]*(-25))+$signed(in_buffer[1]*(-6))+$signed(in_buffer[2]*(-30))+$signed(in_buffer[3]*(-27))+$signed(in_buffer[4]*(11))+$signed(in_buffer[5]*(7))+$signed(in_buffer[6]*(12))+$signed(in_buffer[7]*(-18))+$signed(in_buffer[8]*(-3))+$signed(in_buffer[9]*(-6))+$signed(in_buffer[10]*(14))+$signed(in_buffer[11]*(15))+$signed(in_buffer[12]*(-29))+$signed(in_buffer[13]*(-29))+$signed(in_buffer[14]*(10))+$signed(in_buffer[15]*(-27))+$signed(in_buffer[16]*(2))+$signed(in_buffer[17]*(-7))+$signed(in_buffer[18]*(-17))+$signed(in_buffer[19]*(3))+$signed(in_buffer[20]*(-2))+$signed(in_buffer[21]*(7))+$signed(in_buffer[22]*(19))+$signed(in_buffer[23]*(-12))+$signed(in_buffer[24]*(17));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight55;
assign in_buffer_weight55=$signed(in_buffer[0]*(-6))+$signed(in_buffer[1]*(33))+$signed(in_buffer[2]*(-33))+$signed(in_buffer[3]*(0))+$signed(in_buffer[4]*(12))+$signed(in_buffer[5]*(44))+$signed(in_buffer[6]*(44))+$signed(in_buffer[7]*(62))+$signed(in_buffer[8]*(3))+$signed(in_buffer[9]*(7))+$signed(in_buffer[10]*(-96))+$signed(in_buffer[11]*(-57))+$signed(in_buffer[12]*(-17))+$signed(in_buffer[13]*(0))+$signed(in_buffer[14]*(0))+$signed(in_buffer[15]*(-36))+$signed(in_buffer[16]*(-54))+$signed(in_buffer[17]*(19))+$signed(in_buffer[18]*(-5))+$signed(in_buffer[19]*(-9))+$signed(in_buffer[20]*(101))+$signed(in_buffer[21]*(20))+$signed(in_buffer[22]*(-16))+$signed(in_buffer[23]*(11))+$signed(in_buffer[24]*(32));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight56;
assign in_buffer_weight56=$signed(in_buffer[0]*(-49))+$signed(in_buffer[1]*(33))+$signed(in_buffer[2]*(33))+$signed(in_buffer[3]*(5))+$signed(in_buffer[4]*(-7))+$signed(in_buffer[5]*(-14))+$signed(in_buffer[6]*(18))+$signed(in_buffer[7]*(-32))+$signed(in_buffer[8]*(-15))+$signed(in_buffer[9]*(-7))+$signed(in_buffer[10]*(4))+$signed(in_buffer[11]*(-18))+$signed(in_buffer[12]*(53))+$signed(in_buffer[13]*(65))+$signed(in_buffer[14]*(-17))+$signed(in_buffer[15]*(0))+$signed(in_buffer[16]*(-35))+$signed(in_buffer[17]*(33))+$signed(in_buffer[18]*(10))+$signed(in_buffer[19]*(-55))+$signed(in_buffer[20]*(40))+$signed(in_buffer[21]*(-42))+$signed(in_buffer[22]*(-21))+$signed(in_buffer[23]*(4))+$signed(in_buffer[24]*(106));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight57;
assign in_buffer_weight57=$signed(in_buffer[0]*(-223))+$signed(in_buffer[1]*(-62))+$signed(in_buffer[2]*(18))+$signed(in_buffer[3]*(-5))+$signed(in_buffer[4]*(66))+$signed(in_buffer[5]*(-121))+$signed(in_buffer[6]*(9))+$signed(in_buffer[7]*(32))+$signed(in_buffer[8]*(-37))+$signed(in_buffer[9]*(17))+$signed(in_buffer[10]*(20))+$signed(in_buffer[11]*(-27))+$signed(in_buffer[12]*(70))+$signed(in_buffer[13]*(-16))+$signed(in_buffer[14]*(-144))+$signed(in_buffer[15]*(13))+$signed(in_buffer[16]*(31))+$signed(in_buffer[17]*(-6))+$signed(in_buffer[18]*(-52))+$signed(in_buffer[19]*(52))+$signed(in_buffer[20]*(-20))+$signed(in_buffer[21]*(-26))+$signed(in_buffer[22]*(-21))+$signed(in_buffer[23]*(103))+$signed(in_buffer[24]*(19));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight58;
assign in_buffer_weight58=$signed(in_buffer[0]*(-47))+$signed(in_buffer[1]*(-12))+$signed(in_buffer[2]*(10))+$signed(in_buffer[3]*(25))+$signed(in_buffer[4]*(7))+$signed(in_buffer[5]*(-45))+$signed(in_buffer[6]*(60))+$signed(in_buffer[7]*(9))+$signed(in_buffer[8]*(-39))+$signed(in_buffer[9]*(0))+$signed(in_buffer[10]*(25))+$signed(in_buffer[11]*(54))+$signed(in_buffer[12]*(-106))+$signed(in_buffer[13]*(21))+$signed(in_buffer[14]*(-32))+$signed(in_buffer[15]*(-4))+$signed(in_buffer[16]*(-18))+$signed(in_buffer[17]*(-75))+$signed(in_buffer[18]*(24))+$signed(in_buffer[19]*(12))+$signed(in_buffer[20]*(-53))+$signed(in_buffer[21]*(39))+$signed(in_buffer[22]*(75))+$signed(in_buffer[23]*(12))+$signed(in_buffer[24]*(24));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight59;
assign in_buffer_weight59=$signed(in_buffer[0]*(71))+$signed(in_buffer[1]*(93))+$signed(in_buffer[2]*(0))+$signed(in_buffer[3]*(8))+$signed(in_buffer[4]*(7))+$signed(in_buffer[5]*(-80))+$signed(in_buffer[6]*(-67))+$signed(in_buffer[7]*(-18))+$signed(in_buffer[8]*(-7))+$signed(in_buffer[9]*(-3))+$signed(in_buffer[10]*(-18))+$signed(in_buffer[11]*(15))+$signed(in_buffer[12]*(97))+$signed(in_buffer[13]*(-66))+$signed(in_buffer[14]*(41))+$signed(in_buffer[15]*(58))+$signed(in_buffer[16]*(32))+$signed(in_buffer[17]*(-15))+$signed(in_buffer[18]*(41))+$signed(in_buffer[19]*(29))+$signed(in_buffer[20]*(-50))+$signed(in_buffer[21]*(-22))+$signed(in_buffer[22]*(-13))+$signed(in_buffer[23]*(-53))+$signed(in_buffer[24]*(-86));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight60;
assign in_buffer_weight60=$signed(in_buffer[0]*(-32))+$signed(in_buffer[1]*(6))+$signed(in_buffer[2]*(33))+$signed(in_buffer[3]*(-19))+$signed(in_buffer[4]*(-53))+$signed(in_buffer[5]*(16))+$signed(in_buffer[6]*(-28))+$signed(in_buffer[7]*(-3))+$signed(in_buffer[8]*(6))+$signed(in_buffer[9]*(-34))+$signed(in_buffer[10]*(25))+$signed(in_buffer[11]*(-46))+$signed(in_buffer[12]*(53))+$signed(in_buffer[13]*(-30))+$signed(in_buffer[14]*(-27))+$signed(in_buffer[15]*(1))+$signed(in_buffer[16]*(28))+$signed(in_buffer[17]*(-9))+$signed(in_buffer[18]*(38))+$signed(in_buffer[19]*(38))+$signed(in_buffer[20]*(-1))+$signed(in_buffer[21]*(13))+$signed(in_buffer[22]*(28))+$signed(in_buffer[23]*(8))+$signed(in_buffer[24]*(-1));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight61;
assign in_buffer_weight61=$signed(in_buffer[0]*(-24))+$signed(in_buffer[1]*(12))+$signed(in_buffer[2]*(26))+$signed(in_buffer[3]*(35))+$signed(in_buffer[4]*(-13))+$signed(in_buffer[5]*(19))+$signed(in_buffer[6]*(-9))+$signed(in_buffer[7]*(-32))+$signed(in_buffer[8]*(-44))+$signed(in_buffer[9]*(-24))+$signed(in_buffer[10]*(14))+$signed(in_buffer[11]*(32))+$signed(in_buffer[12]*(-31))+$signed(in_buffer[13]*(18))+$signed(in_buffer[14]*(88))+$signed(in_buffer[15]*(-13))+$signed(in_buffer[16]*(49))+$signed(in_buffer[17]*(9))+$signed(in_buffer[18]*(-25))+$signed(in_buffer[19]*(1))+$signed(in_buffer[20]*(51))+$signed(in_buffer[21]*(28))+$signed(in_buffer[22]*(-46))+$signed(in_buffer[23]*(-20))+$signed(in_buffer[24]*(31));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight62;
assign in_buffer_weight62=$signed(in_buffer[0]*(7))+$signed(in_buffer[1]*(-14))+$signed(in_buffer[2]*(4))+$signed(in_buffer[3]*(-25))+$signed(in_buffer[4]*(20))+$signed(in_buffer[5]*(-20))+$signed(in_buffer[6]*(25))+$signed(in_buffer[7]*(-26))+$signed(in_buffer[8]*(20))+$signed(in_buffer[9]*(27))+$signed(in_buffer[10]*(8))+$signed(in_buffer[11]*(-24))+$signed(in_buffer[12]*(-17))+$signed(in_buffer[13]*(-9))+$signed(in_buffer[14]*(-16))+$signed(in_buffer[15]*(-10))+$signed(in_buffer[16]*(-22))+$signed(in_buffer[17]*(3))+$signed(in_buffer[18]*(-14))+$signed(in_buffer[19]*(12))+$signed(in_buffer[20]*(3))+$signed(in_buffer[21]*(0))+$signed(in_buffer[22]*(11))+$signed(in_buffer[23]*(-4))+$signed(in_buffer[24]*(16));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight63;
assign in_buffer_weight63=$signed(in_buffer[0]*(69))+$signed(in_buffer[1]*(26))+$signed(in_buffer[2]*(-34))+$signed(in_buffer[3]*(20))+$signed(in_buffer[4]*(10))+$signed(in_buffer[5]*(-8))+$signed(in_buffer[6]*(37))+$signed(in_buffer[7]*(-53))+$signed(in_buffer[8]*(-1))+$signed(in_buffer[9]*(-7))+$signed(in_buffer[10]*(18))+$signed(in_buffer[11]*(-5))+$signed(in_buffer[12]*(32))+$signed(in_buffer[13]*(70))+$signed(in_buffer[14]*(-20))+$signed(in_buffer[15]*(-4))+$signed(in_buffer[16]*(0))+$signed(in_buffer[17]*(27))+$signed(in_buffer[18]*(-21))+$signed(in_buffer[19]*(-102))+$signed(in_buffer[20]*(-8))+$signed(in_buffer[21]*(-25))+$signed(in_buffer[22]*(15))+$signed(in_buffer[23]*(-26))+$signed(in_buffer[24]*(2));
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
wire signed [DATA_WIDTH-1:0]   weight_bias10;
wire signed [DATA_WIDTH-1:0]   weight_bias11;
wire signed [DATA_WIDTH-1:0]   weight_bias12;
wire signed [DATA_WIDTH-1:0]   weight_bias13;
wire signed [DATA_WIDTH-1:0]   weight_bias14;
wire signed [DATA_WIDTH-1:0]   weight_bias15;
wire signed [DATA_WIDTH-1:0]   weight_bias16;
wire signed [DATA_WIDTH-1:0]   weight_bias17;
wire signed [DATA_WIDTH-1:0]   weight_bias18;
wire signed [DATA_WIDTH-1:0]   weight_bias19;
wire signed [DATA_WIDTH-1:0]   weight_bias20;
wire signed [DATA_WIDTH-1:0]   weight_bias21;
wire signed [DATA_WIDTH-1:0]   weight_bias22;
wire signed [DATA_WIDTH-1:0]   weight_bias23;
wire signed [DATA_WIDTH-1:0]   weight_bias24;
wire signed [DATA_WIDTH-1:0]   weight_bias25;
wire signed [DATA_WIDTH-1:0]   weight_bias26;
wire signed [DATA_WIDTH-1:0]   weight_bias27;
wire signed [DATA_WIDTH-1:0]   weight_bias28;
wire signed [DATA_WIDTH-1:0]   weight_bias29;
wire signed [DATA_WIDTH-1:0]   weight_bias30;
wire signed [DATA_WIDTH-1:0]   weight_bias31;
wire signed [DATA_WIDTH-1:0]   weight_bias32;
wire signed [DATA_WIDTH-1:0]   weight_bias33;
wire signed [DATA_WIDTH-1:0]   weight_bias34;
wire signed [DATA_WIDTH-1:0]   weight_bias35;
wire signed [DATA_WIDTH-1:0]   weight_bias36;
wire signed [DATA_WIDTH-1:0]   weight_bias37;
wire signed [DATA_WIDTH-1:0]   weight_bias38;
wire signed [DATA_WIDTH-1:0]   weight_bias39;
wire signed [DATA_WIDTH-1:0]   weight_bias40;
wire signed [DATA_WIDTH-1:0]   weight_bias41;
wire signed [DATA_WIDTH-1:0]   weight_bias42;
wire signed [DATA_WIDTH-1:0]   weight_bias43;
wire signed [DATA_WIDTH-1:0]   weight_bias44;
wire signed [DATA_WIDTH-1:0]   weight_bias45;
wire signed [DATA_WIDTH-1:0]   weight_bias46;
wire signed [DATA_WIDTH-1:0]   weight_bias47;
wire signed [DATA_WIDTH-1:0]   weight_bias48;
wire signed [DATA_WIDTH-1:0]   weight_bias49;
wire signed [DATA_WIDTH-1:0]   weight_bias50;
wire signed [DATA_WIDTH-1:0]   weight_bias51;
wire signed [DATA_WIDTH-1:0]   weight_bias52;
wire signed [DATA_WIDTH-1:0]   weight_bias53;
wire signed [DATA_WIDTH-1:0]   weight_bias54;
wire signed [DATA_WIDTH-1:0]   weight_bias55;
wire signed [DATA_WIDTH-1:0]   weight_bias56;
wire signed [DATA_WIDTH-1:0]   weight_bias57;
wire signed [DATA_WIDTH-1:0]   weight_bias58;
wire signed [DATA_WIDTH-1:0]   weight_bias59;
wire signed [DATA_WIDTH-1:0]   weight_bias60;
wire signed [DATA_WIDTH-1:0]   weight_bias61;
wire signed [DATA_WIDTH-1:0]   weight_bias62;
wire signed [DATA_WIDTH-1:0]   weight_bias63;
assign weight_bias0=in_buffer_weight0+(-17);
assign weight_bias1=in_buffer_weight1+(-39);
assign weight_bias2=in_buffer_weight2+(16);
assign weight_bias3=in_buffer_weight3+(29);
assign weight_bias4=in_buffer_weight4+(-34);
assign weight_bias5=in_buffer_weight5+(27);
assign weight_bias6=in_buffer_weight6+(11);
assign weight_bias7=in_buffer_weight7+(-31);
assign weight_bias8=in_buffer_weight8+(47);
assign weight_bias9=in_buffer_weight9+(44);
assign weight_bias10=in_buffer_weight10+(5);
assign weight_bias11=in_buffer_weight11+(24);
assign weight_bias12=in_buffer_weight12+(67);
assign weight_bias13=in_buffer_weight13+(13);
assign weight_bias14=in_buffer_weight14+(44);
assign weight_bias15=in_buffer_weight15+(51);
assign weight_bias16=in_buffer_weight16+(-6);
assign weight_bias17=in_buffer_weight17+(38);
assign weight_bias18=in_buffer_weight18+(41);
assign weight_bias19=in_buffer_weight19+(-27);
assign weight_bias20=in_buffer_weight20+(-21);
assign weight_bias21=in_buffer_weight21+(15);
assign weight_bias22=in_buffer_weight22+(-20);
assign weight_bias23=in_buffer_weight23+(7);
assign weight_bias24=in_buffer_weight24+(-57);
assign weight_bias25=in_buffer_weight25+(-12);
assign weight_bias26=in_buffer_weight26+(69);
assign weight_bias27=in_buffer_weight27+(4);
assign weight_bias28=in_buffer_weight28+(-5);
assign weight_bias29=in_buffer_weight29+(-14);
assign weight_bias30=in_buffer_weight30+(34);
assign weight_bias31=in_buffer_weight31+(37);
assign weight_bias32=in_buffer_weight32+(-20);
assign weight_bias33=in_buffer_weight33+(-17);
assign weight_bias34=in_buffer_weight34+(0);
assign weight_bias35=in_buffer_weight35+(-4);
assign weight_bias36=in_buffer_weight36+(8);
assign weight_bias37=in_buffer_weight37+(-28);
assign weight_bias38=in_buffer_weight38+(-58);
assign weight_bias39=in_buffer_weight39+(-16);
assign weight_bias40=in_buffer_weight40+(-11);
assign weight_bias41=in_buffer_weight41+(-42);
assign weight_bias42=in_buffer_weight42+(17);
assign weight_bias43=in_buffer_weight43+(-44);
assign weight_bias44=in_buffer_weight44+(73);
assign weight_bias45=in_buffer_weight45+(-5);
assign weight_bias46=in_buffer_weight46+(-5);
assign weight_bias47=in_buffer_weight47+(43);
assign weight_bias48=in_buffer_weight48+(-27);
assign weight_bias49=in_buffer_weight49+(-64);
assign weight_bias50=in_buffer_weight50+(16);
assign weight_bias51=in_buffer_weight51+(-53);
assign weight_bias52=in_buffer_weight52+(-58);
assign weight_bias53=in_buffer_weight53+(-1);
assign weight_bias54=in_buffer_weight54+(-19);
assign weight_bias55=in_buffer_weight55+(94);
assign weight_bias56=in_buffer_weight56+(66);
assign weight_bias57=in_buffer_weight57+(9);
assign weight_bias58=in_buffer_weight58+(72);
assign weight_bias59=in_buffer_weight59+(-34);
assign weight_bias60=in_buffer_weight60+(4);
assign weight_bias61=in_buffer_weight61+(17);
assign weight_bias62=in_buffer_weight62+(-1);
assign weight_bias63=in_buffer_weight63+(-19);
wire signed [DATA_WIDTH-1:0]   bias_relu0;
wire signed [DATA_WIDTH-1:0]   bias_relu1;
wire signed [DATA_WIDTH-1:0]   bias_relu2;
wire signed [DATA_WIDTH-1:0]   bias_relu3;
wire signed [DATA_WIDTH-1:0]   bias_relu4;
wire signed [DATA_WIDTH-1:0]   bias_relu5;
wire signed [DATA_WIDTH-1:0]   bias_relu6;
wire signed [DATA_WIDTH-1:0]   bias_relu7;
wire signed [DATA_WIDTH-1:0]   bias_relu8;
wire signed [DATA_WIDTH-1:0]   bias_relu9;
wire signed [DATA_WIDTH-1:0]   bias_relu10;
wire signed [DATA_WIDTH-1:0]   bias_relu11;
wire signed [DATA_WIDTH-1:0]   bias_relu12;
wire signed [DATA_WIDTH-1:0]   bias_relu13;
wire signed [DATA_WIDTH-1:0]   bias_relu14;
wire signed [DATA_WIDTH-1:0]   bias_relu15;
wire signed [DATA_WIDTH-1:0]   bias_relu16;
wire signed [DATA_WIDTH-1:0]   bias_relu17;
wire signed [DATA_WIDTH-1:0]   bias_relu18;
wire signed [DATA_WIDTH-1:0]   bias_relu19;
wire signed [DATA_WIDTH-1:0]   bias_relu20;
wire signed [DATA_WIDTH-1:0]   bias_relu21;
wire signed [DATA_WIDTH-1:0]   bias_relu22;
wire signed [DATA_WIDTH-1:0]   bias_relu23;
wire signed [DATA_WIDTH-1:0]   bias_relu24;
wire signed [DATA_WIDTH-1:0]   bias_relu25;
wire signed [DATA_WIDTH-1:0]   bias_relu26;
wire signed [DATA_WIDTH-1:0]   bias_relu27;
wire signed [DATA_WIDTH-1:0]   bias_relu28;
wire signed [DATA_WIDTH-1:0]   bias_relu29;
wire signed [DATA_WIDTH-1:0]   bias_relu30;
wire signed [DATA_WIDTH-1:0]   bias_relu31;
wire signed [DATA_WIDTH-1:0]   bias_relu32;
wire signed [DATA_WIDTH-1:0]   bias_relu33;
wire signed [DATA_WIDTH-1:0]   bias_relu34;
wire signed [DATA_WIDTH-1:0]   bias_relu35;
wire signed [DATA_WIDTH-1:0]   bias_relu36;
wire signed [DATA_WIDTH-1:0]   bias_relu37;
wire signed [DATA_WIDTH-1:0]   bias_relu38;
wire signed [DATA_WIDTH-1:0]   bias_relu39;
wire signed [DATA_WIDTH-1:0]   bias_relu40;
wire signed [DATA_WIDTH-1:0]   bias_relu41;
wire signed [DATA_WIDTH-1:0]   bias_relu42;
wire signed [DATA_WIDTH-1:0]   bias_relu43;
wire signed [DATA_WIDTH-1:0]   bias_relu44;
wire signed [DATA_WIDTH-1:0]   bias_relu45;
wire signed [DATA_WIDTH-1:0]   bias_relu46;
wire signed [DATA_WIDTH-1:0]   bias_relu47;
wire signed [DATA_WIDTH-1:0]   bias_relu48;
wire signed [DATA_WIDTH-1:0]   bias_relu49;
wire signed [DATA_WIDTH-1:0]   bias_relu50;
wire signed [DATA_WIDTH-1:0]   bias_relu51;
wire signed [DATA_WIDTH-1:0]   bias_relu52;
wire signed [DATA_WIDTH-1:0]   bias_relu53;
wire signed [DATA_WIDTH-1:0]   bias_relu54;
wire signed [DATA_WIDTH-1:0]   bias_relu55;
wire signed [DATA_WIDTH-1:0]   bias_relu56;
wire signed [DATA_WIDTH-1:0]   bias_relu57;
wire signed [DATA_WIDTH-1:0]   bias_relu58;
wire signed [DATA_WIDTH-1:0]   bias_relu59;
wire signed [DATA_WIDTH-1:0]   bias_relu60;
wire signed [DATA_WIDTH-1:0]   bias_relu61;
wire signed [DATA_WIDTH-1:0]   bias_relu62;
wire signed [DATA_WIDTH-1:0]   bias_relu63;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign bias_relu32=(weight_bias32[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias32;
assign bias_relu33=(weight_bias33[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias33;
assign bias_relu34=(weight_bias34[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias34;
assign bias_relu35=(weight_bias35[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias35;
assign bias_relu36=(weight_bias36[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias36;
assign bias_relu37=(weight_bias37[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias37;
assign bias_relu38=(weight_bias38[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias38;
assign bias_relu39=(weight_bias39[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias39;
assign bias_relu40=(weight_bias40[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias40;
assign bias_relu41=(weight_bias41[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias41;
assign bias_relu42=(weight_bias42[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias42;
assign bias_relu43=(weight_bias43[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias43;
assign bias_relu44=(weight_bias44[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias44;
assign bias_relu45=(weight_bias45[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias45;
assign bias_relu46=(weight_bias46[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias46;
assign bias_relu47=(weight_bias47[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias47;
assign bias_relu48=(weight_bias48[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias48;
assign bias_relu49=(weight_bias49[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias49;
assign bias_relu50=(weight_bias50[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias50;
assign bias_relu51=(weight_bias51[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias51;
assign bias_relu52=(weight_bias52[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias52;
assign bias_relu53=(weight_bias53[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias53;
assign bias_relu54=(weight_bias54[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias54;
assign bias_relu55=(weight_bias55[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias55;
assign bias_relu56=(weight_bias56[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias56;
assign bias_relu57=(weight_bias57[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias57;
assign bias_relu58=(weight_bias58[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias58;
assign bias_relu59=(weight_bias59[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias59;
assign bias_relu60=(weight_bias60[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias60;
assign bias_relu61=(weight_bias61[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias61;
assign bias_relu62=(weight_bias62[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias62;
assign bias_relu63=(weight_bias63[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias63;
assign layer_out={bias_relu63,bias_relu62,bias_relu61,bias_relu60,bias_relu59,bias_relu58,bias_relu57,bias_relu56,bias_relu55,bias_relu54,bias_relu53,bias_relu52,bias_relu51,bias_relu50,bias_relu49,bias_relu48,bias_relu47,bias_relu46,bias_relu45,bias_relu44,bias_relu43,bias_relu42,bias_relu41,bias_relu40,bias_relu39,bias_relu38,bias_relu37,bias_relu36,bias_relu35,bias_relu34,bias_relu33,bias_relu32,bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule