module layer1_tcbcnn_121_25x64x10
(
    input clk,
    input rst,
    input [1728-1:0] layer_in,
    input valid,
    output  reg ready,
    output [36*10-1:0] layer_out
);
parameter DATA_WIDTH = 36;
parameter INPUT_DATA_CNT   =   64;
reg    signed [27-1:0]  in_buffer[0:INPUT_DATA_CNT-1];
genvar j;
generate
for(j=0;j<INPUT_DATA_CNT;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=layer_in[j*27+26:j*27+0];
                    end
            end
    end
endgenerate
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0$signed(in_buffer[0]*(10));$signed(in_buffer[1]*(42));$signed(in_buffer[2]*(8));$signed(in_buffer[3]*(-2));$signed(in_buffer[4]*(-24));$signed(in_buffer[5]*(-5));$signed(in_buffer[6]*(-6));$signed(in_buffer[7]*(-28));$signed(in_buffer[8]*(-146));$signed(in_buffer[9]*(-20));$signed(in_buffer[10]*(-38));$signed(in_buffer[11]*(27));$signed(in_buffer[12]*(-110));$signed(in_buffer[13]*(45));$signed(in_buffer[14]*(95));$signed(in_buffer[15]*(-161));$signed(in_buffer[16]*(23));$signed(in_buffer[17]*(7));$signed(in_buffer[18]*(-60));$signed(in_buffer[19]*(-74));$signed(in_buffer[20]*(8));$signed(in_buffer[21]*(-166));$signed(in_buffer[22]*(-21));$signed(in_buffer[23]*(-43));$signed(in_buffer[24]*(-62));$signed(in_buffer[25]*(58));$signed(in_buffer[26]*(2));$signed(in_buffer[27]*(0));$signed(in_buffer[28]*(-76));$signed(in_buffer[29]*(33));$signed(in_buffer[30]*(21));$signed(in_buffer[31]*(22));$signed(in_buffer[32]*(-41));$signed(in_buffer[33]*(31));$signed(in_buffer[34]*(-55));$signed(in_buffer[35]*(-108));$signed(in_buffer[36]*(10));$signed(in_buffer[37]*(53));$signed(in_buffer[38]*(0));$signed(in_buffer[39]*(-12));$signed(in_buffer[40]*(9));$signed(in_buffer[41]*(55));$signed(in_buffer[42]*(43));$signed(in_buffer[43]*(115));$signed(in_buffer[44]*(41));$signed(in_buffer[45]*(-16));$signed(in_buffer[46]*(34));$signed(in_buffer[47]*(-14));$signed(in_buffer[48]*(-113));$signed(in_buffer[49]*(27));$signed(in_buffer[50]*(0));$signed(in_buffer[51]*(-46));$signed(in_buffer[52]*(53));$signed(in_buffer[53]*(-7));$signed(in_buffer[54]*(5));$signed(in_buffer[55]*(20));$signed(in_buffer[56]*(38));$signed(in_buffer[57]*(3));$signed(in_buffer[58]*(-63));$signed(in_buffer[59]*(-24));$signed(in_buffer[60]*(-86));$signed(in_buffer[61]*(-55));$signed(in_buffer[62]*(-27));$signed(in_buffer[63]*(12));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0$signed(in_buffer[0]*(-7));$signed(in_buffer[1]*(-29));$signed(in_buffer[2]*(-51));$signed(in_buffer[3]*(0));$signed(in_buffer[4]*(35));$signed(in_buffer[5]*(-12));$signed(in_buffer[6]*(-17));$signed(in_buffer[7]*(101));$signed(in_buffer[8]*(-55));$signed(in_buffer[9]*(10));$signed(in_buffer[10]*(0));$signed(in_buffer[11]*(75));$signed(in_buffer[12]*(144));$signed(in_buffer[13]*(-17));$signed(in_buffer[14]*(75));$signed(in_buffer[15]*(-22));$signed(in_buffer[16]*(71));$signed(in_buffer[17]*(11));$signed(in_buffer[18]*(57));$signed(in_buffer[19]*(-34));$signed(in_buffer[20]*(-104));$signed(in_buffer[21]*(-7));$signed(in_buffer[22]*(24));$signed(in_buffer[23]*(-115));$signed(in_buffer[24]*(18));$signed(in_buffer[25]*(101));$signed(in_buffer[26]*(-9));$signed(in_buffer[27]*(-42));$signed(in_buffer[28]*(56));$signed(in_buffer[29]*(-16));$signed(in_buffer[30]*(-38));$signed(in_buffer[31]*(-26));$signed(in_buffer[32]*(-101));$signed(in_buffer[33]*(-77));$signed(in_buffer[34]*(-124));$signed(in_buffer[35]*(-106));$signed(in_buffer[36]*(-10));$signed(in_buffer[37]*(7));$signed(in_buffer[38]*(-10));$signed(in_buffer[39]*(-38));$signed(in_buffer[40]*(-24));$signed(in_buffer[41]*(-17));$signed(in_buffer[42]*(-54));$signed(in_buffer[43]*(9));$signed(in_buffer[44]*(19));$signed(in_buffer[45]*(48));$signed(in_buffer[46]*(-42));$signed(in_buffer[47]*(-145));$signed(in_buffer[48]*(76));$signed(in_buffer[49]*(63));$signed(in_buffer[50]*(92));$signed(in_buffer[51]*(59));$signed(in_buffer[52]*(-31));$signed(in_buffer[53]*(11));$signed(in_buffer[54]*(-106));$signed(in_buffer[55]*(-110));$signed(in_buffer[56]*(-7));$signed(in_buffer[57]*(5));$signed(in_buffer[58]*(47));$signed(in_buffer[59]*(-71));$signed(in_buffer[60]*(93));$signed(in_buffer[61]*(-19));$signed(in_buffer[62]*(24));$signed(in_buffer[63]*(-15));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0$signed(in_buffer[0]*(-3));$signed(in_buffer[1]*(-2));$signed(in_buffer[2]*(21));$signed(in_buffer[3]*(-21));$signed(in_buffer[4]*(-45));$signed(in_buffer[5]*(-6));$signed(in_buffer[6]*(38));$signed(in_buffer[7]*(-56));$signed(in_buffer[8]*(47));$signed(in_buffer[9]*(92));$signed(in_buffer[10]*(-31));$signed(in_buffer[11]*(-12));$signed(in_buffer[12]*(-72));$signed(in_buffer[13]*(-34));$signed(in_buffer[14]*(-61));$signed(in_buffer[15]*(-75));$signed(in_buffer[16]*(5));$signed(in_buffer[17]*(18));$signed(in_buffer[18]*(74));$signed(in_buffer[19]*(-62));$signed(in_buffer[20]*(-36));$signed(in_buffer[21]*(41));$signed(in_buffer[22]*(8));$signed(in_buffer[23]*(20));$signed(in_buffer[24]*(15));$signed(in_buffer[25]*(28));$signed(in_buffer[26]*(16));$signed(in_buffer[27]*(7));$signed(in_buffer[28]*(24));$signed(in_buffer[29]*(1));$signed(in_buffer[30]*(32));$signed(in_buffer[31]*(-43));$signed(in_buffer[32]*(1));$signed(in_buffer[33]*(-36));$signed(in_buffer[34]*(133));$signed(in_buffer[35]*(-21));$signed(in_buffer[36]*(-11));$signed(in_buffer[37]*(10));$signed(in_buffer[38]*(-9));$signed(in_buffer[39]*(-26));$signed(in_buffer[40]*(10));$signed(in_buffer[41]*(18));$signed(in_buffer[42]*(11));$signed(in_buffer[43]*(-23));$signed(in_buffer[44]*(16));$signed(in_buffer[45]*(-42));$signed(in_buffer[46]*(-5));$signed(in_buffer[47]*(92));$signed(in_buffer[48]*(-84));$signed(in_buffer[49]*(5));$signed(in_buffer[50]*(32));$signed(in_buffer[51]*(3));$signed(in_buffer[52]*(14));$signed(in_buffer[53]*(-12));$signed(in_buffer[54]*(-15));$signed(in_buffer[55]*(14));$signed(in_buffer[56]*(31));$signed(in_buffer[57]*(-8));$signed(in_buffer[58]*(12));$signed(in_buffer[59]*(4));$signed(in_buffer[60]*(-103));$signed(in_buffer[61]*(37));$signed(in_buffer[62]*(21));$signed(in_buffer[63]*(-123));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0$signed(in_buffer[0]*(-7));$signed(in_buffer[1]*(-44));$signed(in_buffer[2]*(16));$signed(in_buffer[3]*(-71));$signed(in_buffer[4]*(-40));$signed(in_buffer[5]*(8));$signed(in_buffer[6]*(-21));$signed(in_buffer[7]*(-62));$signed(in_buffer[8]*(40));$signed(in_buffer[9]*(-53));$signed(in_buffer[10]*(-34));$signed(in_buffer[11]*(-24));$signed(in_buffer[12]*(-62));$signed(in_buffer[13]*(68));$signed(in_buffer[14]*(-124));$signed(in_buffer[15]*(40));$signed(in_buffer[16]*(5));$signed(in_buffer[17]*(-15));$signed(in_buffer[18]*(83));$signed(in_buffer[19]*(56));$signed(in_buffer[20]*(0));$signed(in_buffer[21]*(69));$signed(in_buffer[22]*(-12));$signed(in_buffer[23]*(24));$signed(in_buffer[24]*(59));$signed(in_buffer[25]*(16));$signed(in_buffer[26]*(6));$signed(in_buffer[27]*(4));$signed(in_buffer[28]*(-23));$signed(in_buffer[29]*(-4));$signed(in_buffer[30]*(-15));$signed(in_buffer[31]*(-75));$signed(in_buffer[32]*(-17));$signed(in_buffer[33]*(-14));$signed(in_buffer[34]*(-1));$signed(in_buffer[35]*(30));$signed(in_buffer[36]*(-3));$signed(in_buffer[37]*(39));$signed(in_buffer[38]*(-27));$signed(in_buffer[39]*(-65));$signed(in_buffer[40]*(16));$signed(in_buffer[41]*(57));$signed(in_buffer[42]*(36));$signed(in_buffer[43]*(-51));$signed(in_buffer[44]*(-87));$signed(in_buffer[45]*(19));$signed(in_buffer[46]*(36));$signed(in_buffer[47]*(23));$signed(in_buffer[48]*(6));$signed(in_buffer[49]*(6));$signed(in_buffer[50]*(-36));$signed(in_buffer[51]*(47));$signed(in_buffer[52]*(-8));$signed(in_buffer[53]*(-2));$signed(in_buffer[54]*(2));$signed(in_buffer[55]*(-31));$signed(in_buffer[56]*(-28));$signed(in_buffer[57]*(2));$signed(in_buffer[58]*(13));$signed(in_buffer[59]*(-5));$signed(in_buffer[60]*(-69));$signed(in_buffer[61]*(32));$signed(in_buffer[62]*(22));$signed(in_buffer[63]*(-60));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0$signed(in_buffer[0]*(-2));$signed(in_buffer[1]*(26));$signed(in_buffer[2]*(-55));$signed(in_buffer[3]*(-23));$signed(in_buffer[4]*(30));$signed(in_buffer[5]*(-8));$signed(in_buffer[6]*(27));$signed(in_buffer[7]*(-193));$signed(in_buffer[8]*(54));$signed(in_buffer[9]*(32));$signed(in_buffer[10]*(33));$signed(in_buffer[11]*(61));$signed(in_buffer[12]*(32));$signed(in_buffer[13]*(-30));$signed(in_buffer[14]*(19));$signed(in_buffer[15]*(61));$signed(in_buffer[16]*(-97));$signed(in_buffer[17]*(-41));$signed(in_buffer[18]*(-242));$signed(in_buffer[19]*(28));$signed(in_buffer[20]*(14));$signed(in_buffer[21]*(-26));$signed(in_buffer[22]*(-33));$signed(in_buffer[23]*(7));$signed(in_buffer[24]*(-93));$signed(in_buffer[25]*(-23));$signed(in_buffer[26]*(2));$signed(in_buffer[27]*(-59));$signed(in_buffer[28]*(27));$signed(in_buffer[29]*(1));$signed(in_buffer[30]*(-29));$signed(in_buffer[31]*(-68));$signed(in_buffer[32]*(-4));$signed(in_buffer[33]*(29));$signed(in_buffer[34]*(-65));$signed(in_buffer[35]*(38));$signed(in_buffer[36]*(-9));$signed(in_buffer[37]*(-19));$signed(in_buffer[38]*(0));$signed(in_buffer[39]*(41));$signed(in_buffer[40]*(-32));$signed(in_buffer[41]*(-24));$signed(in_buffer[42]*(-2));$signed(in_buffer[43]*(-35));$signed(in_buffer[44]*(54));$signed(in_buffer[45]*(-58));$signed(in_buffer[46]*(-38));$signed(in_buffer[47]*(44));$signed(in_buffer[48]*(119));$signed(in_buffer[49]*(7));$signed(in_buffer[50]*(7));$signed(in_buffer[51]*(-21));$signed(in_buffer[52]*(-69));$signed(in_buffer[53]*(-2));$signed(in_buffer[54]*(-60));$signed(in_buffer[55]*(-40));$signed(in_buffer[56]*(-6));$signed(in_buffer[57]*(6));$signed(in_buffer[58]*(29));$signed(in_buffer[59]*(84));$signed(in_buffer[60]*(-2));$signed(in_buffer[61]*(-93));$signed(in_buffer[62]*(-1));$signed(in_buffer[63]*(-74));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0$signed(in_buffer[0]*(-13));$signed(in_buffer[1]*(36));$signed(in_buffer[2]*(-49));$signed(in_buffer[3]*(0));$signed(in_buffer[4]*(15));$signed(in_buffer[5]*(-12));$signed(in_buffer[6]*(-34));$signed(in_buffer[7]*(160));$signed(in_buffer[8]*(22));$signed(in_buffer[9]*(-79));$signed(in_buffer[10]*(-40));$signed(in_buffer[11]*(-88));$signed(in_buffer[12]*(59));$signed(in_buffer[13]*(28));$signed(in_buffer[14]*(-34));$signed(in_buffer[15]*(29));$signed(in_buffer[16]*(54));$signed(in_buffer[17]*(30));$signed(in_buffer[18]*(-71));$signed(in_buffer[19]*(53));$signed(in_buffer[20]*(-10));$signed(in_buffer[21]*(45));$signed(in_buffer[22]*(-11));$signed(in_buffer[23]*(25));$signed(in_buffer[24]*(-32));$signed(in_buffer[25]*(6));$signed(in_buffer[26]*(-1));$signed(in_buffer[27]*(-65));$signed(in_buffer[28]*(25));$signed(in_buffer[29]*(0));$signed(in_buffer[30]*(-40));$signed(in_buffer[31]*(44));$signed(in_buffer[32]*(-4));$signed(in_buffer[33]*(-21));$signed(in_buffer[34]*(48));$signed(in_buffer[35]*(-8));$signed(in_buffer[36]*(-5));$signed(in_buffer[37]*(29));$signed(in_buffer[38]*(-20));$signed(in_buffer[39]*(12));$signed(in_buffer[40]*(-2));$signed(in_buffer[41]*(-7));$signed(in_buffer[42]*(35));$signed(in_buffer[43]*(-177));$signed(in_buffer[44]*(0));$signed(in_buffer[45]*(15));$signed(in_buffer[46]*(54));$signed(in_buffer[47]*(10));$signed(in_buffer[48]*(-47));$signed(in_buffer[49]*(-79));$signed(in_buffer[50]*(42));$signed(in_buffer[51]*(2));$signed(in_buffer[52]*(13));$signed(in_buffer[53]*(13));$signed(in_buffer[54]*(43));$signed(in_buffer[55]*(23));$signed(in_buffer[56]*(-12));$signed(in_buffer[57]*(5));$signed(in_buffer[58]*(13));$signed(in_buffer[59]*(-14));$signed(in_buffer[60]*(92));$signed(in_buffer[61]*(28));$signed(in_buffer[62]*(-65));$signed(in_buffer[63]*(40));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0$signed(in_buffer[0]*(9));$signed(in_buffer[1]*(-8));$signed(in_buffer[2]*(31));$signed(in_buffer[3]*(10));$signed(in_buffer[4]*(39));$signed(in_buffer[5]*(-13));$signed(in_buffer[6]*(26));$signed(in_buffer[7]*(41));$signed(in_buffer[8]*(-39));$signed(in_buffer[9]*(63));$signed(in_buffer[10]*(35));$signed(in_buffer[11]*(0));$signed(in_buffer[12]*(84));$signed(in_buffer[13]*(-23));$signed(in_buffer[14]*(82));$signed(in_buffer[15]*(-139));$signed(in_buffer[16]*(-16));$signed(in_buffer[17]*(-160));$signed(in_buffer[18]*(-174));$signed(in_buffer[19]*(-72));$signed(in_buffer[20]*(0));$signed(in_buffer[21]*(-153));$signed(in_buffer[22]*(38));$signed(in_buffer[23]*(-170));$signed(in_buffer[24]*(-81));$signed(in_buffer[25]*(-1));$signed(in_buffer[26]*(0));$signed(in_buffer[27]*(-79));$signed(in_buffer[28]*(56));$signed(in_buffer[29]*(34));$signed(in_buffer[30]*(20));$signed(in_buffer[31]*(25));$signed(in_buffer[32]*(17));$signed(in_buffer[33]*(34));$signed(in_buffer[34]*(60));$signed(in_buffer[35]*(-9));$signed(in_buffer[36]*(5));$signed(in_buffer[37]*(-70));$signed(in_buffer[38]*(-2));$signed(in_buffer[39]*(40));$signed(in_buffer[40]*(-33));$signed(in_buffer[41]*(-24));$signed(in_buffer[42]*(-63));$signed(in_buffer[43]*(-10));$signed(in_buffer[44]*(-14));$signed(in_buffer[45]*(-52));$signed(in_buffer[46]*(-41));$signed(in_buffer[47]*(18));$signed(in_buffer[48]*(4));$signed(in_buffer[49]*(-3));$signed(in_buffer[50]*(-150));$signed(in_buffer[51]*(-3));$signed(in_buffer[52]*(24));$signed(in_buffer[53]*(-3));$signed(in_buffer[54]*(20));$signed(in_buffer[55]*(-7));$signed(in_buffer[56]*(-6));$signed(in_buffer[57]*(5));$signed(in_buffer[58]*(-36));$signed(in_buffer[59]*(33));$signed(in_buffer[60]*(41));$signed(in_buffer[61]*(-39));$signed(in_buffer[62]*(-166));$signed(in_buffer[63]*(168));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0$signed(in_buffer[0]*(13));$signed(in_buffer[1]*(-26));$signed(in_buffer[2]*(-35));$signed(in_buffer[3]*(38));$signed(in_buffer[4]*(-12));$signed(in_buffer[5]*(-4));$signed(in_buffer[6]*(-51));$signed(in_buffer[7]*(-19));$signed(in_buffer[8]*(-5));$signed(in_buffer[9]*(-36));$signed(in_buffer[10]*(-25));$signed(in_buffer[11]*(8));$signed(in_buffer[12]*(-162));$signed(in_buffer[13]*(-8));$signed(in_buffer[14]*(6));$signed(in_buffer[15]*(21));$signed(in_buffer[16]*(-2));$signed(in_buffer[17]*(32));$signed(in_buffer[18]*(87));$signed(in_buffer[19]*(-43));$signed(in_buffer[20]*(33));$signed(in_buffer[21]*(77));$signed(in_buffer[22]*(44));$signed(in_buffer[23]*(50));$signed(in_buffer[24]*(-4));$signed(in_buffer[25]*(67));$signed(in_buffer[26]*(11));$signed(in_buffer[27]*(39));$signed(in_buffer[28]*(66));$signed(in_buffer[29]*(-44));$signed(in_buffer[30]*(-3));$signed(in_buffer[31]*(92));$signed(in_buffer[32]*(-90));$signed(in_buffer[33]*(50));$signed(in_buffer[34]*(30));$signed(in_buffer[35]*(14));$signed(in_buffer[36]*(1));$signed(in_buffer[37]*(30));$signed(in_buffer[38]*(1));$signed(in_buffer[39]*(1));$signed(in_buffer[40]*(14));$signed(in_buffer[41]*(8));$signed(in_buffer[42]*(-14));$signed(in_buffer[43]*(61));$signed(in_buffer[44]*(43));$signed(in_buffer[45]*(7));$signed(in_buffer[46]*(-67));$signed(in_buffer[47]*(3));$signed(in_buffer[48]*(-10));$signed(in_buffer[49]*(-91));$signed(in_buffer[50]*(-33));$signed(in_buffer[51]*(-47));$signed(in_buffer[52]*(-5));$signed(in_buffer[53]*(7));$signed(in_buffer[54]*(71));$signed(in_buffer[55]*(-27));$signed(in_buffer[56]*(-70));$signed(in_buffer[57]*(-1));$signed(in_buffer[58]*(-23));$signed(in_buffer[59]*(-82));$signed(in_buffer[60]*(-117));$signed(in_buffer[61]*(-89));$signed(in_buffer[62]*(29));$signed(in_buffer[63]*(-80));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0$signed(in_buffer[0]*(9));$signed(in_buffer[1]*(0));$signed(in_buffer[2]*(24));$signed(in_buffer[3]*(13));$signed(in_buffer[4]*(10));$signed(in_buffer[5]*(13));$signed(in_buffer[6]*(-52));$signed(in_buffer[7]*(-33));$signed(in_buffer[8]*(-45));$signed(in_buffer[9]*(-54));$signed(in_buffer[10]*(21));$signed(in_buffer[11]*(-64));$signed(in_buffer[12]*(-42));$signed(in_buffer[13]*(-61));$signed(in_buffer[14]*(-42));$signed(in_buffer[15]*(-12));$signed(in_buffer[16]*(8));$signed(in_buffer[17]*(16));$signed(in_buffer[18]*(-19));$signed(in_buffer[19]*(44));$signed(in_buffer[20]*(11));$signed(in_buffer[21]*(-14));$signed(in_buffer[22]*(-5));$signed(in_buffer[23]*(-8));$signed(in_buffer[24]*(47));$signed(in_buffer[25]*(-92));$signed(in_buffer[26]*(14));$signed(in_buffer[27]*(36));$signed(in_buffer[28]*(-17));$signed(in_buffer[29]*(42));$signed(in_buffer[30]*(29));$signed(in_buffer[31]*(-1));$signed(in_buffer[32]*(79));$signed(in_buffer[33]*(-2));$signed(in_buffer[34]*(-26));$signed(in_buffer[35]*(-9));$signed(in_buffer[36]*(-1));$signed(in_buffer[37]*(-74));$signed(in_buffer[38]*(-22));$signed(in_buffer[39]*(-10));$signed(in_buffer[40]*(29));$signed(in_buffer[41]*(-87));$signed(in_buffer[42]*(18));$signed(in_buffer[43]*(0));$signed(in_buffer[44]*(-76));$signed(in_buffer[45]*(31));$signed(in_buffer[46]*(25));$signed(in_buffer[47]*(-88));$signed(in_buffer[48]*(-83));$signed(in_buffer[49]*(8));$signed(in_buffer[50]*(-72));$signed(in_buffer[51]*(16));$signed(in_buffer[52]*(7));$signed(in_buffer[53]*(-12));$signed(in_buffer[54]*(-48));$signed(in_buffer[55]*(8));$signed(in_buffer[56]*(-9));$signed(in_buffer[57]*(2));$signed(in_buffer[58]*(37));$signed(in_buffer[59]*(-101));$signed(in_buffer[60]*(-39));$signed(in_buffer[61]*(60));$signed(in_buffer[62]*(-17));$signed(in_buffer[63]*(-8));;
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0$signed(in_buffer[0]*(-15));$signed(in_buffer[1]*(-4));$signed(in_buffer[2]*(-6));$signed(in_buffer[3]*(33));$signed(in_buffer[4]*(-1));$signed(in_buffer[5]*(1));$signed(in_buffer[6]*(-77));$signed(in_buffer[7]*(-43));$signed(in_buffer[8]*(0));$signed(in_buffer[9]*(37));$signed(in_buffer[10]*(12));$signed(in_buffer[11]*(79));$signed(in_buffer[12]*(-163));$signed(in_buffer[13]*(-20));$signed(in_buffer[14]*(3));$signed(in_buffer[15]*(42));$signed(in_buffer[16]*(-7));$signed(in_buffer[17]*(17));$signed(in_buffer[18]*(-95));$signed(in_buffer[19]*(-64));$signed(in_buffer[20]*(24));$signed(in_buffer[21]*(-78));$signed(in_buffer[22]*(-133));$signed(in_buffer[23]*(36));$signed(in_buffer[24]*(30));$signed(in_buffer[25]*(-194));$signed(in_buffer[26]*(11));$signed(in_buffer[27]*(50));$signed(in_buffer[28]*(-215));$signed(in_buffer[29]*(-72));$signed(in_buffer[30]*(4));$signed(in_buffer[31]*(-78));$signed(in_buffer[32]*(-27));$signed(in_buffer[33]*(24));$signed(in_buffer[34]*(-200));$signed(in_buffer[35]*(40));$signed(in_buffer[36]*(-17));$signed(in_buffer[37]*(-20));$signed(in_buffer[38]*(-2));$signed(in_buffer[39]*(6));$signed(in_buffer[40]*(1));$signed(in_buffer[41]*(-3));$signed(in_buffer[42]*(-24));$signed(in_buffer[43]*(56));$signed(in_buffer[44]*(31));$signed(in_buffer[45]*(3));$signed(in_buffer[46]*(-8));$signed(in_buffer[47]*(-43));$signed(in_buffer[48]*(30));$signed(in_buffer[49]*(42));$signed(in_buffer[50]*(23));$signed(in_buffer[51]*(-37));$signed(in_buffer[52]*(-52));$signed(in_buffer[53]*(-3));$signed(in_buffer[54]*(8));$signed(in_buffer[55]*(4));$signed(in_buffer[56]*(14));$signed(in_buffer[57]*(10));$signed(in_buffer[58]*(11));$signed(in_buffer[59]*(40));$signed(in_buffer[60]*(17));$signed(in_buffer[61]*(-23));$signed(in_buffer[62]*(47));$signed(in_buffer[63]*(-2));;
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias0=in_buffer_weight0+(-9);
assign weight_bias1=in_buffer_weight1+(12);
assign weight_bias2=in_buffer_weight2+(-37);
assign weight_bias3=in_buffer_weight3+(-13);
assign weight_bias4=in_buffer_weight4+(2);
assign weight_bias5=in_buffer_weight5+(19);
assign weight_bias6=in_buffer_weight6+(-11);
assign weight_bias7=in_buffer_weight7+(10);
assign weight_bias8=in_buffer_weight8+(-11);
assign weight_bias9=in_buffer_weight9+(16);
assign layer_out={weight_bias9,weight_bias8,weight_bias7,weight_bias6,weight_bias5,weight_bias4,weight_bias3,weight_bias2,weight_bias1,weight_bias0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule