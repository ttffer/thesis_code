`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/22/2022 05:59:06 PM
// Design Name: 
// Module Name: n13sys5x5_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module n13sys5x5_testbench(

    );
    reg [5:0] word0,word1,word2,word3,word4,word5,word6,word7,word8,word9,word10,word11,word12,word13,word14,word15,word16,word17,word18,word19,word20,word21,word22,word23,word24;
    wire [2:0] d_word0,d_word1,d_word2,d_word3,d_word4,d_word5,d_word6,d_word7,d_word8,d_word9,d_word10,d_word11,d_word12,d_word13,d_word14,d_word15,d_word16,d_word17,d_word18,d_word19,d_word20,d_word21,d_word22,d_word23,d_word24;
    n13sys_5x5 DUT_n13(.IN0(word0),.IN1(word1),.IN2(word2),.IN3(word3),.IN4(word4),.IN5(word5),.IN6(word6),.IN7(word7),.IN8(word8),.IN9(word9),.IN10(word10),.IN11(word11),.IN12(word12),.IN13(word13),.IN14(word14),.IN15(word15),.IN16(word16),.IN17(word17),.IN18(word18),.IN19(word19),.IN20(word20),.IN21(word21),.IN22(word22),.IN23(word23),.IN24(word24),.OUT0(d_word0),.OUT1(d_word1),.OUT2(d_word2),.OUT3(d_word3),.OUT4(d_word4),.OUT5(d_word5),.OUT6(d_word6),.OUT7(d_word7),.OUT8(d_word8),.OUT9(d_word9),.OUT10(d_word10),.OUT11(d_word11),.OUT12(d_word12),.OUT13(d_word13),.OUT14(d_word14),.OUT15(d_word15),.OUT16(d_word16),.OUT17(d_word17),.OUT18(d_word18),.OUT19(d_word19),.OUT20(d_word20),.OUT21(d_word21),.OUT22(d_word22),.OUT23(d_word23),.OUT24(d_word24));
    
    initial begin  
    word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d1;
#10 word0='d6;
 #10 word0='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d1;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d2;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d4;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d8;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d16;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d32;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d12;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d15;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d9;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d5;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d29;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d45;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d27;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d24;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d30;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d18;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d10;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d58;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d38;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d37;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d35;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d47;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d55;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d7;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d53;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d54;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d48;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d60;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d36;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word0='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word1='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word2='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word3='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word4='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word5='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word6='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word7='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word8='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word9='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word10='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word11='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word12='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word13='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word14='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word15='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word16='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word17='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word18='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word19='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word20='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word21='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word22='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word23='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
#10 word24='d20;
#10 word0=6'd0;word1=6'd0;word2=6'd0;word3=6'd0;word4=6'd0;word5=6'd0;word6=6'd0;word7=6'd0;word8=6'd0;word9=6'd0;word10=6'd0;word11=6'd0;word12=6'd0;word13=6'd0;word14=6'd0;word15=6'd0;word16=6'd0;word17=6'd0;word18=6'd0;word19=6'd0;word20=6'd0;word21=6'd0;word22=6'd0;word23=6'd0;word24=6'd0;
  
    $stop;
    end
    
    
endmodule
