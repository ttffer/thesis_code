module layer2_tcb_121x16x10
(
    input clk,
    input rst,
   input valid,
   output  reg ready,
    input [27*16-1:0]  layer_in,
    output [42*10-1:0]   layer_out
);
parameter DATA_WIDTH   =   42;
reg [DATA_WIDTH-1:0]    layer_in_buffer    [0:16-1];
integer i;
always@(posedge clk )
    begin
        if(rst)
            begin
                for(i=0;i<16;i=i+1)
                    begin
                        layer_in_buffer[i]<=0;
                    end
            end
        else
        begin
       layer_in_buffer[0]<=layer_in[26:0];
       layer_in_buffer[1]<=layer_in[53:27];
       layer_in_buffer[2]<=layer_in[80:54];
       layer_in_buffer[3]<=layer_in[107:81];
       layer_in_buffer[4]<=layer_in[134:108];
       layer_in_buffer[5]<=layer_in[161:135];
       layer_in_buffer[6]<=layer_in[188:162];
       layer_in_buffer[7]<=layer_in[215:189];
       layer_in_buffer[8]<=layer_in[242:216];
       layer_in_buffer[9]<=layer_in[269:243];
       layer_in_buffer[10]<=layer_in[296:270];
       layer_in_buffer[11]<=layer_in[323:297];
       layer_in_buffer[12]<=layer_in[350:324];
       layer_in_buffer[13]<=layer_in[377:351];
       layer_in_buffer[14]<=layer_in[404:378];
       layer_in_buffer[15]<=layer_in[431:405];
        end
   end

wire [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0-(0+(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<3)-(layer_in_buffer[0]<<7)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<12)+(layer_in_buffer[0]<<13))-(0-(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<4)+(layer_in_buffer[1]<<7)+(layer_in_buffer[1]<<11))+(0+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<5)-(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<11))-(0+(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<5)+(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<11)+(layer_in_buffer[3]<<13))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<9))+(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<1)-(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<10))+(0-(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<11))-(0-(layer_in_buffer[7]<<1)+(layer_in_buffer[7]<<6)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<9))+(0+(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<9)+(layer_in_buffer[8]<<12))+(0-(layer_in_buffer[9]<<0)+(layer_in_buffer[9]<<5)-(layer_in_buffer[9]<<8)-(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<12)+(layer_in_buffer[9]<<13))+(0+(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<4)-(layer_in_buffer[10]<<6)+(layer_in_buffer[10]<<9)+(layer_in_buffer[10]<<12))-(0+(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<2)-(layer_in_buffer[11]<<4)-(layer_in_buffer[11]<<7)+(layer_in_buffer[11]<<11))-(0+(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<13))+(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<11))-(0-(layer_in_buffer[14]<<1)+(layer_in_buffer[14]<<6)+(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<9))-(0+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<5)+(layer_in_buffer[15]<<9)+(layer_in_buffer[15]<<12));
wire [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0-(0+(layer_in_buffer[0]<<5)-(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<13))+(0+(layer_in_buffer[1]<<1)+(layer_in_buffer[1]<<4)+(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<13))+(0+(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<11))-(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<1)+(layer_in_buffer[3]<<5)-(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<12)+(layer_in_buffer[3]<<14))+(0+(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<11))+(0+(layer_in_buffer[5]<<6)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<10)+(layer_in_buffer[5]<<12))-(0+(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<12)+(layer_in_buffer[6]<<14))-(0+(layer_in_buffer[7]<<0)-(layer_in_buffer[7]<<2)-(layer_in_buffer[7]<<4)-(layer_in_buffer[7]<<6)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<12)+(layer_in_buffer[7]<<14))+(0-(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<2)-(layer_in_buffer[8]<<4)+(layer_in_buffer[8]<<7)-(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<12)+(layer_in_buffer[8]<<13))-(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6)-(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<11)+(layer_in_buffer[9]<<13))-(0+(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<1)-(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<8)-(layer_in_buffer[10]<<11)+(layer_in_buffer[10]<<14))-(0+(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<14))+(0+(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<5)+(layer_in_buffer[12]<<7)+(layer_in_buffer[12]<<8)+(layer_in_buffer[12]<<11)+(layer_in_buffer[12]<<12))+(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<2)-(layer_in_buffer[13]<<4)-(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<11))-(0+(layer_in_buffer[14]<<3)+(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<7)+(layer_in_buffer[14]<<9))+(0+(layer_in_buffer[15]<<1)-(layer_in_buffer[15]<<3)-(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<9)+(layer_in_buffer[15]<<11));
wire [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0-(0-(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)-(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<9))+(0+(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<6)+(layer_in_buffer[1]<<9)+(layer_in_buffer[1]<<11))-(0+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<3)+(layer_in_buffer[2]<<5)-(layer_in_buffer[2]<<7)+(layer_in_buffer[2]<<10)+(layer_in_buffer[2]<<13))+(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<4)-(layer_in_buffer[3]<<7)+(layer_in_buffer[3]<<10))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<3)+(layer_in_buffer[4]<<6)+(layer_in_buffer[4]<<10))+(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<5)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<10)+(layer_in_buffer[5]<<11))-(0+(layer_in_buffer[6]<<0)-(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<5)+(layer_in_buffer[6]<<7)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<12))-(0+(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<11))+(0-(layer_in_buffer[8]<<1)+(layer_in_buffer[8]<<4)+(layer_in_buffer[8]<<5)+(layer_in_buffer[8]<<8)-(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<13))-(0-(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<4)+(layer_in_buffer[9]<<6)-(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<14))-(0+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7))+(0+(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<6)-(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<12))-(0+(layer_in_buffer[12]<<1)+(layer_in_buffer[12]<<6)+(layer_in_buffer[12]<<9)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<13))-(0-(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<5)+(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<8))-(0-(layer_in_buffer[14]<<1)-(layer_in_buffer[14]<<3)-(layer_in_buffer[14]<<5)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<10))-(0+(layer_in_buffer[15]<<3)-(layer_in_buffer[15]<<5)-(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<11)+(layer_in_buffer[15]<<13));
wire [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0-(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<4)-(layer_in_buffer[0]<<9)+(layer_in_buffer[0]<<12))-(0+(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<10)+(layer_in_buffer[1]<<13))+(0+(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<12))-(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6)+(layer_in_buffer[3]<<9))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<9))+(0+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<7)-(layer_in_buffer[5]<<10)+(layer_in_buffer[5]<<13))+(0-(layer_in_buffer[6]<<0)-(layer_in_buffer[6]<<2)-(layer_in_buffer[6]<<4)-(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<12))-(0+(layer_in_buffer[7]<<0)-(layer_in_buffer[7]<<4)-(layer_in_buffer[7]<<6)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<13))+(0-(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<7)+(layer_in_buffer[8]<<9)+(layer_in_buffer[8]<<10))-(0+(layer_in_buffer[9]<<5)+(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<11)+(layer_in_buffer[9]<<14))-(0+(layer_in_buffer[10]<<3)+(layer_in_buffer[10]<<4)-(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<12)+(layer_in_buffer[10]<<13))+(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<7)+(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<12))+(0+(layer_in_buffer[12]<<6)+(layer_in_buffer[12]<<7)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<12))+(0-(layer_in_buffer[13]<<0)-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<5)+(layer_in_buffer[13]<<11))+(0+(layer_in_buffer[14]<<1)-(layer_in_buffer[14]<<3)-(layer_in_buffer[14]<<6)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<11))-(0-(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<5)-(layer_in_buffer[15]<<9)+(layer_in_buffer[15]<<13));
wire [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0-(0+(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<2)-(layer_in_buffer[0]<<4)-(layer_in_buffer[0]<<7)+(layer_in_buffer[0]<<11))+(0-(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<6)+(layer_in_buffer[1]<<12))+(0+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<2)-(layer_in_buffer[2]<<5)-(layer_in_buffer[2]<<7)-(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<11)+(layer_in_buffer[2]<<12))+(0+(layer_in_buffer[3]<<1)-(layer_in_buffer[3]<<5)-(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<13))-(0-(layer_in_buffer[4]<<1)-(layer_in_buffer[4]<<3)-(layer_in_buffer[4]<<5)+(layer_in_buffer[4]<<9)+(layer_in_buffer[4]<<10))+(0-(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<10))-(0+(layer_in_buffer[6]<<1)+(layer_in_buffer[6]<<2)-(layer_in_buffer[6]<<5)-(layer_in_buffer[6]<<7)-(layer_in_buffer[6]<<9)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<12))+(0+(layer_in_buffer[7]<<0)-(layer_in_buffer[7]<<4)-(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<12))+(0-(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<6)-(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<11))-(0+(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<5)-(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<12)+(layer_in_buffer[9]<<14))+(0+(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)-(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<8)+(layer_in_buffer[10]<<10))-(0-(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<5)-(layer_in_buffer[11]<<7)-(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<12))+(0+(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<4)+(layer_in_buffer[12]<<6)+(layer_in_buffer[12]<<11)+(layer_in_buffer[12]<<12))+(0+(layer_in_buffer[13]<<4)+(layer_in_buffer[13]<<5)+(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<10))-(0-(layer_in_buffer[14]<<1)-(layer_in_buffer[14]<<3)-(layer_in_buffer[14]<<5)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<10))-(0+(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<11)+(layer_in_buffer[15]<<14));
wire [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0+(0+(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<8)-(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<13)+(layer_in_buffer[0]<<14))-(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<3)-(layer_in_buffer[1]<<6)-(layer_in_buffer[1]<<9)+(layer_in_buffer[1]<<12)+(layer_in_buffer[1]<<13))-(0-(layer_in_buffer[2]<<2)-(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<12))+(0+(layer_in_buffer[3]<<1)+(layer_in_buffer[3]<<2)-(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<11))-(0+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<5)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<10))-(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<8)-(layer_in_buffer[5]<<10)+(layer_in_buffer[5]<<13)+(layer_in_buffer[5]<<14))-(0-(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<11))-(0-(layer_in_buffer[7]<<1)+(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<4)+(layer_in_buffer[7]<<7)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<11)+(layer_in_buffer[7]<<12))+(0+(layer_in_buffer[8]<<0)-(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<5)+(layer_in_buffer[8]<<6)-(layer_in_buffer[8]<<9)+(layer_in_buffer[8]<<12)+(layer_in_buffer[8]<<13))+(0+(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<6)-(layer_in_buffer[9]<<9)+(layer_in_buffer[9]<<12))+(0+(layer_in_buffer[10]<<1)-(layer_in_buffer[10]<<5)-(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<13))+(0-(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<10)+(layer_in_buffer[11]<<12)+(layer_in_buffer[11]<<13))+(0-(layer_in_buffer[12]<<2)-(layer_in_buffer[12]<<4)+(layer_in_buffer[12]<<7)+(layer_in_buffer[12]<<13))+(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<9))+(0+(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<6)+(layer_in_buffer[14]<<7)+(layer_in_buffer[14]<<11))+(0+(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<2)-(layer_in_buffer[15]<<5)-(layer_in_buffer[15]<<7)-(layer_in_buffer[15]<<9)+(layer_in_buffer[15]<<11)+(layer_in_buffer[15]<<12));
wire [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0-(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)-(layer_in_buffer[0]<<4)-(layer_in_buffer[0]<<6)+(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<9)+(layer_in_buffer[0]<<12)+(layer_in_buffer[0]<<14))+(0+(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<7)-(layer_in_buffer[1]<<10)+(layer_in_buffer[1]<<13))-(0+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<3)-(layer_in_buffer[2]<<5)-(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<12))-(0+(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<7)+(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<12)+(layer_in_buffer[3]<<13))+(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<9))+(0+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<9))+(0-(layer_in_buffer[6]<<2)-(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<7)+(layer_in_buffer[6]<<13))+(0-(layer_in_buffer[7]<<2)-(layer_in_buffer[7]<<5)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<12))-(0+(layer_in_buffer[8]<<1)-(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<6)-(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<11)+(layer_in_buffer[8]<<12))+(0-(layer_in_buffer[9]<<1)-(layer_in_buffer[9]<<3)-(layer_in_buffer[9]<<5)-(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<12)+(layer_in_buffer[9]<<13))+(0-(layer_in_buffer[10]<<1)-(layer_in_buffer[10]<<3)-(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<9)+(layer_in_buffer[10]<<10))+(0+(layer_in_buffer[11]<<1)-(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<9))+(0-(layer_in_buffer[12]<<1)+(layer_in_buffer[12]<<4)+(layer_in_buffer[12]<<5)+(layer_in_buffer[12]<<8)-(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<13))-(0+(layer_in_buffer[13]<<2)-(layer_in_buffer[13]<<5)+(layer_in_buffer[13]<<10))+(0+(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<5)+(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<10))-(0-(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<4)+(layer_in_buffer[15]<<5)+(layer_in_buffer[15]<<8)-(layer_in_buffer[15]<<10)+(layer_in_buffer[15]<<13));
wire [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0-(0-(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<7)+(layer_in_buffer[0]<<9)+(layer_in_buffer[0]<<12))-(0+(layer_in_buffer[1]<<0)+(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<5)-(layer_in_buffer[1]<<9)-(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<14))+(0-(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<4)-(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<9)+(layer_in_buffer[2]<<12))+(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<1)-(layer_in_buffer[3]<<4)-(layer_in_buffer[3]<<6)-(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<11))-(0+(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<3)+(layer_in_buffer[4]<<8))-(0+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<6)-(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<12))+(0+(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<6)-(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<14))+(0+(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<4)+(layer_in_buffer[7]<<6)+(layer_in_buffer[7]<<11)+(layer_in_buffer[7]<<12))-(0+(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<1)-(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<6)-(layer_in_buffer[8]<<9)+(layer_in_buffer[8]<<13)+(layer_in_buffer[8]<<14))-(0+(layer_in_buffer[9]<<2)-(layer_in_buffer[9]<<4)+(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<9)-(layer_in_buffer[9]<<13)+(layer_in_buffer[9]<<16))-(0+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<2)-(layer_in_buffer[10]<<6)+(layer_in_buffer[10]<<13))-(0-(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<4)-(layer_in_buffer[11]<<6)-(layer_in_buffer[11]<<8)-(layer_in_buffer[11]<<10)+(layer_in_buffer[11]<<14))-(0-(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<3)-(layer_in_buffer[12]<<6)-(layer_in_buffer[12]<<8)-(layer_in_buffer[12]<<11)+(layer_in_buffer[12]<<14))-(0+(layer_in_buffer[13]<<3)-(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<11))+(0+(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<3)+(layer_in_buffer[14]<<5)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<10))+(0-(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<5)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<9)+(layer_in_buffer[15]<<13));
wire [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0+(0+(layer_in_buffer[0]<<1)-(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<12)+(layer_in_buffer[0]<<14))-(0+(layer_in_buffer[1]<<1)+(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<7))+(0+(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<7)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<11)+(layer_in_buffer[2]<<12))+(0+(layer_in_buffer[3]<<5)+(layer_in_buffer[3]<<6)+(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<11))+(0-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<9)+(layer_in_buffer[4]<<10))+(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<11))-(0+(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<2)-(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<12)+(layer_in_buffer[6]<<13))+(0-(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<10)+(layer_in_buffer[7]<<11))-(0+(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<1)+(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<9)+(layer_in_buffer[8]<<11)+(layer_in_buffer[8]<<13))-(0+(layer_in_buffer[9]<<0)+(layer_in_buffer[9]<<3)+(layer_in_buffer[9]<<6)+(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<13))-(0+(layer_in_buffer[10]<<3)-(layer_in_buffer[10]<<6)+(layer_in_buffer[10]<<11))+(0+(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<1)-(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<12))-(0-(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<8)+(layer_in_buffer[12]<<13)+(layer_in_buffer[12]<<14))+(0+(layer_in_buffer[13]<<1)-(layer_in_buffer[13]<<3)-(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<9)+(layer_in_buffer[13]<<11))+(0+(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<1)+(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<6))-(0+(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<3)-(layer_in_buffer[15]<<5)-(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<12));
wire [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0-(0+(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<1)-(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<7)+(layer_in_buffer[0]<<9)-(layer_in_buffer[0]<<12)+(layer_in_buffer[0]<<15))-(0-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<7)-(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<15))-(0+(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<3)-(layer_in_buffer[2]<<7)+(layer_in_buffer[2]<<10)+(layer_in_buffer[2]<<13)+(layer_in_buffer[2]<<14))+(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6)+(layer_in_buffer[3]<<9))+(0+(layer_in_buffer[4]<<3)+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<9))+(0+(layer_in_buffer[5]<<1)+(layer_in_buffer[5]<<5)-(layer_in_buffer[5]<<8)+(layer_in_buffer[5]<<11))-(0+(layer_in_buffer[6]<<1)+(layer_in_buffer[6]<<4)-(layer_in_buffer[6]<<6)-(layer_in_buffer[6]<<9)-(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<14))+(0-(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<13))-(0+(layer_in_buffer[8]<<3)+(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<12)+(layer_in_buffer[8]<<13))-(0+(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<4)+(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<13))+(0+(layer_in_buffer[10]<<0)+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<13))-(0-(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<6)-(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<11)+(layer_in_buffer[11]<<12))+(0+(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<13))+(0+(layer_in_buffer[13]<<3)-(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<11))-(0+(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<1)-(layer_in_buffer[14]<<7)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<10))+(0+(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<4)+(layer_in_buffer[15]<<10)+(layer_in_buffer[15]<<12));
wire [DATA_WIDTH-1:0]   weight_bias0;
assign weight_bias0=in_buffer_weight0+(-581);
wire [DATA_WIDTH-1:0]   weight_bias1;
assign weight_bias1=in_buffer_weight1+(-747);
wire [DATA_WIDTH-1:0]   weight_bias2;
assign weight_bias2=in_buffer_weight2+(2241);
wire [DATA_WIDTH-1:0]   weight_bias3;
assign weight_bias3=in_buffer_weight3+(-1577);
wire [DATA_WIDTH-1:0]   weight_bias4;
assign weight_bias4=in_buffer_weight4+(-6889);
wire [DATA_WIDTH-1:0]   weight_bias5;
assign weight_bias5=in_buffer_weight5+(4565);
wire [DATA_WIDTH-1:0]   weight_bias6;
assign weight_bias6=in_buffer_weight6+(-2490);
wire [DATA_WIDTH-1:0]   weight_bias7;
assign weight_bias7=in_buffer_weight7+(6640);
wire [DATA_WIDTH-1:0]   weight_bias8;
assign weight_bias8=in_buffer_weight8+(-1992);
wire [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias9=in_buffer_weight9+(-5893);
assign layer_out={
            weight_bias9,
            weight_bias8,
            weight_bias7,
            weight_bias6,
            weight_bias5,
            weight_bias4,
            weight_bias3,
            weight_bias2,
            weight_bias1,
            weight_bias0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule
