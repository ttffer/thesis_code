module n29sys(input [13:0]IN0,input [13:0]IN1,output [9:0]OUT0,output [9:0]OUT1,