module con_tcb
    #(
        parameter   OUTPUT_BIT  =   19,
                    OUTPUT_NODE =   100,
                    DATA_WIDTH  =   19,
                    IMG_SZ    =   11*11
)
(
    input   clk,
    input   rst,
    input   [IMG_SZ*8-1:0]   img,
    input   valid,
    output  reg ready,
    output [OUTPUT_BIT*OUTPUT_NODE-1:0] layer_out
);

reg    signed [8-1:0]  in_buffer[0:IMG_SZ-1];
genvar j;
generate
for(j=0;j<IMG_SZ;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=img[j*8+7:j*8+0];
                    end
            end
    end
endgenerate
//wire declatation
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight0;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight1;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight2;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight3;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight4;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight5;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight6;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight7;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight8;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight9;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight10;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight11;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight12;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight13;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight14;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight15;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight16;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight17;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight18;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight19;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight20;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight21;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight22;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight23;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight24;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight25;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight26;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight27;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight28;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight29;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight30;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight31;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight32;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight33;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight34;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight35;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight36;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight37;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight38;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight39;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight40;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight41;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight42;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight43;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight44;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight45;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight46;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight47;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight48;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight49;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight50;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight51;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight52;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight53;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight54;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight55;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight56;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight57;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight58;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight59;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight60;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight61;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight62;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight63;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight64;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight65;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight66;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight67;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight68;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight69;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight70;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight71;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight72;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight73;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight74;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight75;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight76;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight77;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight78;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight79;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight80;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight81;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight82;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight83;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight84;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight85;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight86;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight87;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight88;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight89;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight90;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight91;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight92;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight93;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight94;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight95;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight96;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight97;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight98;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight99;
assign in_buffer_weight0=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<5)+(in_buffer[0]<<8))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<2)+(in_buffer[1]<<8))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<8))+(0+(in_buffer[12]<<2)+(in_buffer[12]<<4)+(in_buffer[12]<<5)+(in_buffer[12]<<8));
assign in_buffer_weight1=0+(0+(in_buffer[1]<<0)+(in_buffer[1]<<3)+(in_buffer[1]<<5)+(in_buffer[1]<<8))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<2)+(in_buffer[2]<<8))+(0-(in_buffer[12]<<0)+(in_buffer[12]<<8))+(0+(in_buffer[13]<<2)+(in_buffer[13]<<4)+(in_buffer[13]<<5)+(in_buffer[13]<<8));
assign in_buffer_weight2=0+(0+(in_buffer[2]<<0)+(in_buffer[2]<<3)+(in_buffer[2]<<5)+(in_buffer[2]<<8))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<2)+(in_buffer[3]<<8))+(0-(in_buffer[13]<<0)+(in_buffer[13]<<8))+(0+(in_buffer[14]<<2)+(in_buffer[14]<<4)+(in_buffer[14]<<5)+(in_buffer[14]<<8));
assign in_buffer_weight3=0+(0+(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<5)+(in_buffer[3]<<8))+(0+(in_buffer[4]<<1)+(in_buffer[4]<<2)+(in_buffer[4]<<8))+(0-(in_buffer[14]<<0)+(in_buffer[14]<<8))+(0+(in_buffer[15]<<2)+(in_buffer[15]<<4)+(in_buffer[15]<<5)+(in_buffer[15]<<8));
assign in_buffer_weight4=0+(0+(in_buffer[4]<<0)+(in_buffer[4]<<3)+(in_buffer[4]<<5)+(in_buffer[4]<<8))+(0+(in_buffer[5]<<1)+(in_buffer[5]<<2)+(in_buffer[5]<<8))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<8))+(0+(in_buffer[16]<<2)+(in_buffer[16]<<4)+(in_buffer[16]<<5)+(in_buffer[16]<<8));
assign in_buffer_weight5=0+(0+(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<5)+(in_buffer[5]<<8))+(0+(in_buffer[6]<<1)+(in_buffer[6]<<2)+(in_buffer[6]<<8))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<8))+(0+(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<5)+(in_buffer[17]<<8));
assign in_buffer_weight6=0+(0+(in_buffer[6]<<0)+(in_buffer[6]<<3)+(in_buffer[6]<<5)+(in_buffer[6]<<8))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<2)+(in_buffer[7]<<8))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<8))+(0+(in_buffer[18]<<2)+(in_buffer[18]<<4)+(in_buffer[18]<<5)+(in_buffer[18]<<8));
assign in_buffer_weight7=0+(0+(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<5)+(in_buffer[7]<<8))+(0+(in_buffer[8]<<1)+(in_buffer[8]<<2)+(in_buffer[8]<<8))+(0-(in_buffer[18]<<0)+(in_buffer[18]<<8))+(0+(in_buffer[19]<<2)+(in_buffer[19]<<4)+(in_buffer[19]<<5)+(in_buffer[19]<<8));
assign in_buffer_weight8=0+(0+(in_buffer[8]<<0)+(in_buffer[8]<<3)+(in_buffer[8]<<5)+(in_buffer[8]<<8))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<2)+(in_buffer[9]<<8))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<8))+(0+(in_buffer[20]<<2)+(in_buffer[20]<<4)+(in_buffer[20]<<5)+(in_buffer[20]<<8));
assign in_buffer_weight9=0+(0+(in_buffer[9]<<0)+(in_buffer[9]<<3)+(in_buffer[9]<<5)+(in_buffer[9]<<8))+(0+(in_buffer[10]<<1)+(in_buffer[10]<<2)+(in_buffer[10]<<8))+(0-(in_buffer[20]<<0)+(in_buffer[20]<<8))+(0+(in_buffer[21]<<2)+(in_buffer[21]<<4)+(in_buffer[21]<<5)+(in_buffer[21]<<8));
assign in_buffer_weight10=0+(0+(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<5)+(in_buffer[11]<<8))+(0+(in_buffer[12]<<1)+(in_buffer[12]<<2)+(in_buffer[12]<<8))+(0-(in_buffer[22]<<0)+(in_buffer[22]<<8))+(0+(in_buffer[23]<<2)+(in_buffer[23]<<4)+(in_buffer[23]<<5)+(in_buffer[23]<<8));
assign in_buffer_weight11=0+(0+(in_buffer[12]<<0)+(in_buffer[12]<<3)+(in_buffer[12]<<5)+(in_buffer[12]<<8))+(0+(in_buffer[13]<<1)+(in_buffer[13]<<2)+(in_buffer[13]<<8))+(0-(in_buffer[23]<<0)+(in_buffer[23]<<8))+(0+(in_buffer[24]<<2)+(in_buffer[24]<<4)+(in_buffer[24]<<5)+(in_buffer[24]<<8));
assign in_buffer_weight12=0+(0+(in_buffer[13]<<0)+(in_buffer[13]<<3)+(in_buffer[13]<<5)+(in_buffer[13]<<8))+(0+(in_buffer[14]<<1)+(in_buffer[14]<<2)+(in_buffer[14]<<8))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<8))+(0+(in_buffer[25]<<2)+(in_buffer[25]<<4)+(in_buffer[25]<<5)+(in_buffer[25]<<8));
assign in_buffer_weight13=0+(0+(in_buffer[14]<<0)+(in_buffer[14]<<3)+(in_buffer[14]<<5)+(in_buffer[14]<<8))+(0+(in_buffer[15]<<1)+(in_buffer[15]<<2)+(in_buffer[15]<<8))+(0-(in_buffer[25]<<0)+(in_buffer[25]<<8))+(0+(in_buffer[26]<<2)+(in_buffer[26]<<4)+(in_buffer[26]<<5)+(in_buffer[26]<<8));
assign in_buffer_weight14=0+(0+(in_buffer[15]<<0)+(in_buffer[15]<<3)+(in_buffer[15]<<5)+(in_buffer[15]<<8))+(0+(in_buffer[16]<<1)+(in_buffer[16]<<2)+(in_buffer[16]<<8))+(0-(in_buffer[26]<<0)+(in_buffer[26]<<8))+(0+(in_buffer[27]<<2)+(in_buffer[27]<<4)+(in_buffer[27]<<5)+(in_buffer[27]<<8));
assign in_buffer_weight15=0+(0+(in_buffer[16]<<0)+(in_buffer[16]<<3)+(in_buffer[16]<<5)+(in_buffer[16]<<8))+(0+(in_buffer[17]<<1)+(in_buffer[17]<<2)+(in_buffer[17]<<8))+(0-(in_buffer[27]<<0)+(in_buffer[27]<<8))+(0+(in_buffer[28]<<2)+(in_buffer[28]<<4)+(in_buffer[28]<<5)+(in_buffer[28]<<8));
assign in_buffer_weight16=0+(0+(in_buffer[17]<<0)+(in_buffer[17]<<3)+(in_buffer[17]<<5)+(in_buffer[17]<<8))+(0+(in_buffer[18]<<1)+(in_buffer[18]<<2)+(in_buffer[18]<<8))+(0-(in_buffer[28]<<0)+(in_buffer[28]<<8))+(0+(in_buffer[29]<<2)+(in_buffer[29]<<4)+(in_buffer[29]<<5)+(in_buffer[29]<<8));
assign in_buffer_weight17=0+(0+(in_buffer[18]<<0)+(in_buffer[18]<<3)+(in_buffer[18]<<5)+(in_buffer[18]<<8))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<2)+(in_buffer[19]<<8))+(0-(in_buffer[29]<<0)+(in_buffer[29]<<8))+(0+(in_buffer[30]<<2)+(in_buffer[30]<<4)+(in_buffer[30]<<5)+(in_buffer[30]<<8));
assign in_buffer_weight18=0+(0+(in_buffer[19]<<0)+(in_buffer[19]<<3)+(in_buffer[19]<<5)+(in_buffer[19]<<8))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<2)+(in_buffer[20]<<8))+(0-(in_buffer[30]<<0)+(in_buffer[30]<<8))+(0+(in_buffer[31]<<2)+(in_buffer[31]<<4)+(in_buffer[31]<<5)+(in_buffer[31]<<8));
assign in_buffer_weight19=0+(0+(in_buffer[20]<<0)+(in_buffer[20]<<3)+(in_buffer[20]<<5)+(in_buffer[20]<<8))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<2)+(in_buffer[21]<<8))+(0-(in_buffer[31]<<0)+(in_buffer[31]<<8))+(0+(in_buffer[32]<<2)+(in_buffer[32]<<4)+(in_buffer[32]<<5)+(in_buffer[32]<<8));
assign in_buffer_weight20=0+(0+(in_buffer[22]<<0)+(in_buffer[22]<<3)+(in_buffer[22]<<5)+(in_buffer[22]<<8))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<2)+(in_buffer[23]<<8))+(0-(in_buffer[33]<<0)+(in_buffer[33]<<8))+(0+(in_buffer[34]<<2)+(in_buffer[34]<<4)+(in_buffer[34]<<5)+(in_buffer[34]<<8));
assign in_buffer_weight21=0+(0+(in_buffer[23]<<0)+(in_buffer[23]<<3)+(in_buffer[23]<<5)+(in_buffer[23]<<8))+(0+(in_buffer[24]<<1)+(in_buffer[24]<<2)+(in_buffer[24]<<8))+(0-(in_buffer[34]<<0)+(in_buffer[34]<<8))+(0+(in_buffer[35]<<2)+(in_buffer[35]<<4)+(in_buffer[35]<<5)+(in_buffer[35]<<8));
assign in_buffer_weight22=0+(0+(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<5)+(in_buffer[24]<<8))+(0+(in_buffer[25]<<1)+(in_buffer[25]<<2)+(in_buffer[25]<<8))+(0-(in_buffer[35]<<0)+(in_buffer[35]<<8))+(0+(in_buffer[36]<<2)+(in_buffer[36]<<4)+(in_buffer[36]<<5)+(in_buffer[36]<<8));
assign in_buffer_weight23=0+(0+(in_buffer[25]<<0)+(in_buffer[25]<<3)+(in_buffer[25]<<5)+(in_buffer[25]<<8))+(0+(in_buffer[26]<<1)+(in_buffer[26]<<2)+(in_buffer[26]<<8))+(0-(in_buffer[36]<<0)+(in_buffer[36]<<8))+(0+(in_buffer[37]<<2)+(in_buffer[37]<<4)+(in_buffer[37]<<5)+(in_buffer[37]<<8));
assign in_buffer_weight24=0+(0+(in_buffer[26]<<0)+(in_buffer[26]<<3)+(in_buffer[26]<<5)+(in_buffer[26]<<8))+(0+(in_buffer[27]<<1)+(in_buffer[27]<<2)+(in_buffer[27]<<8))+(0-(in_buffer[37]<<0)+(in_buffer[37]<<8))+(0+(in_buffer[38]<<2)+(in_buffer[38]<<4)+(in_buffer[38]<<5)+(in_buffer[38]<<8));
assign in_buffer_weight25=0+(0+(in_buffer[27]<<0)+(in_buffer[27]<<3)+(in_buffer[27]<<5)+(in_buffer[27]<<8))+(0+(in_buffer[28]<<1)+(in_buffer[28]<<2)+(in_buffer[28]<<8))+(0-(in_buffer[38]<<0)+(in_buffer[38]<<8))+(0+(in_buffer[39]<<2)+(in_buffer[39]<<4)+(in_buffer[39]<<5)+(in_buffer[39]<<8));
assign in_buffer_weight26=0+(0+(in_buffer[28]<<0)+(in_buffer[28]<<3)+(in_buffer[28]<<5)+(in_buffer[28]<<8))+(0+(in_buffer[29]<<1)+(in_buffer[29]<<2)+(in_buffer[29]<<8))+(0-(in_buffer[39]<<0)+(in_buffer[39]<<8))+(0+(in_buffer[40]<<2)+(in_buffer[40]<<4)+(in_buffer[40]<<5)+(in_buffer[40]<<8));
assign in_buffer_weight27=0+(0+(in_buffer[29]<<0)+(in_buffer[29]<<3)+(in_buffer[29]<<5)+(in_buffer[29]<<8))+(0+(in_buffer[30]<<1)+(in_buffer[30]<<2)+(in_buffer[30]<<8))+(0-(in_buffer[40]<<0)+(in_buffer[40]<<8))+(0+(in_buffer[41]<<2)+(in_buffer[41]<<4)+(in_buffer[41]<<5)+(in_buffer[41]<<8));
assign in_buffer_weight28=0+(0+(in_buffer[30]<<0)+(in_buffer[30]<<3)+(in_buffer[30]<<5)+(in_buffer[30]<<8))+(0+(in_buffer[31]<<1)+(in_buffer[31]<<2)+(in_buffer[31]<<8))+(0-(in_buffer[41]<<0)+(in_buffer[41]<<8))+(0+(in_buffer[42]<<2)+(in_buffer[42]<<4)+(in_buffer[42]<<5)+(in_buffer[42]<<8));
assign in_buffer_weight29=0+(0+(in_buffer[31]<<0)+(in_buffer[31]<<3)+(in_buffer[31]<<5)+(in_buffer[31]<<8))+(0+(in_buffer[32]<<1)+(in_buffer[32]<<2)+(in_buffer[32]<<8))+(0-(in_buffer[42]<<0)+(in_buffer[42]<<8))+(0+(in_buffer[43]<<2)+(in_buffer[43]<<4)+(in_buffer[43]<<5)+(in_buffer[43]<<8));
assign in_buffer_weight30=0+(0+(in_buffer[33]<<0)+(in_buffer[33]<<3)+(in_buffer[33]<<5)+(in_buffer[33]<<8))+(0+(in_buffer[34]<<1)+(in_buffer[34]<<2)+(in_buffer[34]<<8))+(0-(in_buffer[44]<<0)+(in_buffer[44]<<8))+(0+(in_buffer[45]<<2)+(in_buffer[45]<<4)+(in_buffer[45]<<5)+(in_buffer[45]<<8));
assign in_buffer_weight31=0+(0+(in_buffer[34]<<0)+(in_buffer[34]<<3)+(in_buffer[34]<<5)+(in_buffer[34]<<8))+(0+(in_buffer[35]<<1)+(in_buffer[35]<<2)+(in_buffer[35]<<8))+(0-(in_buffer[45]<<0)+(in_buffer[45]<<8))+(0+(in_buffer[46]<<2)+(in_buffer[46]<<4)+(in_buffer[46]<<5)+(in_buffer[46]<<8));
assign in_buffer_weight32=0+(0+(in_buffer[35]<<0)+(in_buffer[35]<<3)+(in_buffer[35]<<5)+(in_buffer[35]<<8))+(0+(in_buffer[36]<<1)+(in_buffer[36]<<2)+(in_buffer[36]<<8))+(0-(in_buffer[46]<<0)+(in_buffer[46]<<8))+(0+(in_buffer[47]<<2)+(in_buffer[47]<<4)+(in_buffer[47]<<5)+(in_buffer[47]<<8));
assign in_buffer_weight33=0+(0+(in_buffer[36]<<0)+(in_buffer[36]<<3)+(in_buffer[36]<<5)+(in_buffer[36]<<8))+(0+(in_buffer[37]<<1)+(in_buffer[37]<<2)+(in_buffer[37]<<8))+(0-(in_buffer[47]<<0)+(in_buffer[47]<<8))+(0+(in_buffer[48]<<2)+(in_buffer[48]<<4)+(in_buffer[48]<<5)+(in_buffer[48]<<8));
assign in_buffer_weight34=0+(0+(in_buffer[37]<<0)+(in_buffer[37]<<3)+(in_buffer[37]<<5)+(in_buffer[37]<<8))+(0+(in_buffer[38]<<1)+(in_buffer[38]<<2)+(in_buffer[38]<<8))+(0-(in_buffer[48]<<0)+(in_buffer[48]<<8))+(0+(in_buffer[49]<<2)+(in_buffer[49]<<4)+(in_buffer[49]<<5)+(in_buffer[49]<<8));
assign in_buffer_weight35=0+(0+(in_buffer[38]<<0)+(in_buffer[38]<<3)+(in_buffer[38]<<5)+(in_buffer[38]<<8))+(0+(in_buffer[39]<<1)+(in_buffer[39]<<2)+(in_buffer[39]<<8))+(0-(in_buffer[49]<<0)+(in_buffer[49]<<8))+(0+(in_buffer[50]<<2)+(in_buffer[50]<<4)+(in_buffer[50]<<5)+(in_buffer[50]<<8));
assign in_buffer_weight36=0+(0+(in_buffer[39]<<0)+(in_buffer[39]<<3)+(in_buffer[39]<<5)+(in_buffer[39]<<8))+(0+(in_buffer[40]<<1)+(in_buffer[40]<<2)+(in_buffer[40]<<8))+(0-(in_buffer[50]<<0)+(in_buffer[50]<<8))+(0+(in_buffer[51]<<2)+(in_buffer[51]<<4)+(in_buffer[51]<<5)+(in_buffer[51]<<8));
assign in_buffer_weight37=0+(0+(in_buffer[40]<<0)+(in_buffer[40]<<3)+(in_buffer[40]<<5)+(in_buffer[40]<<8))+(0+(in_buffer[41]<<1)+(in_buffer[41]<<2)+(in_buffer[41]<<8))+(0-(in_buffer[51]<<0)+(in_buffer[51]<<8))+(0+(in_buffer[52]<<2)+(in_buffer[52]<<4)+(in_buffer[52]<<5)+(in_buffer[52]<<8));
assign in_buffer_weight38=0+(0+(in_buffer[41]<<0)+(in_buffer[41]<<3)+(in_buffer[41]<<5)+(in_buffer[41]<<8))+(0+(in_buffer[42]<<1)+(in_buffer[42]<<2)+(in_buffer[42]<<8))+(0-(in_buffer[52]<<0)+(in_buffer[52]<<8))+(0+(in_buffer[53]<<2)+(in_buffer[53]<<4)+(in_buffer[53]<<5)+(in_buffer[53]<<8));
assign in_buffer_weight39=0+(0+(in_buffer[42]<<0)+(in_buffer[42]<<3)+(in_buffer[42]<<5)+(in_buffer[42]<<8))+(0+(in_buffer[43]<<1)+(in_buffer[43]<<2)+(in_buffer[43]<<8))+(0-(in_buffer[53]<<0)+(in_buffer[53]<<8))+(0+(in_buffer[54]<<2)+(in_buffer[54]<<4)+(in_buffer[54]<<5)+(in_buffer[54]<<8));
assign in_buffer_weight40=0+(0+(in_buffer[44]<<0)+(in_buffer[44]<<3)+(in_buffer[44]<<5)+(in_buffer[44]<<8))+(0+(in_buffer[45]<<1)+(in_buffer[45]<<2)+(in_buffer[45]<<8))+(0-(in_buffer[55]<<0)+(in_buffer[55]<<8))+(0+(in_buffer[56]<<2)+(in_buffer[56]<<4)+(in_buffer[56]<<5)+(in_buffer[56]<<8));
assign in_buffer_weight41=0+(0+(in_buffer[45]<<0)+(in_buffer[45]<<3)+(in_buffer[45]<<5)+(in_buffer[45]<<8))+(0+(in_buffer[46]<<1)+(in_buffer[46]<<2)+(in_buffer[46]<<8))+(0-(in_buffer[56]<<0)+(in_buffer[56]<<8))+(0+(in_buffer[57]<<2)+(in_buffer[57]<<4)+(in_buffer[57]<<5)+(in_buffer[57]<<8));
assign in_buffer_weight42=0+(0+(in_buffer[46]<<0)+(in_buffer[46]<<3)+(in_buffer[46]<<5)+(in_buffer[46]<<8))+(0+(in_buffer[47]<<1)+(in_buffer[47]<<2)+(in_buffer[47]<<8))+(0-(in_buffer[57]<<0)+(in_buffer[57]<<8))+(0+(in_buffer[58]<<2)+(in_buffer[58]<<4)+(in_buffer[58]<<5)+(in_buffer[58]<<8));
assign in_buffer_weight43=0+(0+(in_buffer[47]<<0)+(in_buffer[47]<<3)+(in_buffer[47]<<5)+(in_buffer[47]<<8))+(0+(in_buffer[48]<<1)+(in_buffer[48]<<2)+(in_buffer[48]<<8))+(0-(in_buffer[58]<<0)+(in_buffer[58]<<8))+(0+(in_buffer[59]<<2)+(in_buffer[59]<<4)+(in_buffer[59]<<5)+(in_buffer[59]<<8));
assign in_buffer_weight44=0+(0+(in_buffer[48]<<0)+(in_buffer[48]<<3)+(in_buffer[48]<<5)+(in_buffer[48]<<8))+(0+(in_buffer[49]<<1)+(in_buffer[49]<<2)+(in_buffer[49]<<8))+(0-(in_buffer[59]<<0)+(in_buffer[59]<<8))+(0+(in_buffer[60]<<2)+(in_buffer[60]<<4)+(in_buffer[60]<<5)+(in_buffer[60]<<8));
assign in_buffer_weight45=0+(0+(in_buffer[49]<<0)+(in_buffer[49]<<3)+(in_buffer[49]<<5)+(in_buffer[49]<<8))+(0+(in_buffer[50]<<1)+(in_buffer[50]<<2)+(in_buffer[50]<<8))+(0-(in_buffer[60]<<0)+(in_buffer[60]<<8))+(0+(in_buffer[61]<<2)+(in_buffer[61]<<4)+(in_buffer[61]<<5)+(in_buffer[61]<<8));
assign in_buffer_weight46=0+(0+(in_buffer[50]<<0)+(in_buffer[50]<<3)+(in_buffer[50]<<5)+(in_buffer[50]<<8))+(0+(in_buffer[51]<<1)+(in_buffer[51]<<2)+(in_buffer[51]<<8))+(0-(in_buffer[61]<<0)+(in_buffer[61]<<8))+(0+(in_buffer[62]<<2)+(in_buffer[62]<<4)+(in_buffer[62]<<5)+(in_buffer[62]<<8));
assign in_buffer_weight47=0+(0+(in_buffer[51]<<0)+(in_buffer[51]<<3)+(in_buffer[51]<<5)+(in_buffer[51]<<8))+(0+(in_buffer[52]<<1)+(in_buffer[52]<<2)+(in_buffer[52]<<8))+(0-(in_buffer[62]<<0)+(in_buffer[62]<<8))+(0+(in_buffer[63]<<2)+(in_buffer[63]<<4)+(in_buffer[63]<<5)+(in_buffer[63]<<8));
assign in_buffer_weight48=0+(0+(in_buffer[52]<<0)+(in_buffer[52]<<3)+(in_buffer[52]<<5)+(in_buffer[52]<<8))+(0+(in_buffer[53]<<1)+(in_buffer[53]<<2)+(in_buffer[53]<<8))+(0-(in_buffer[63]<<0)+(in_buffer[63]<<8))+(0+(in_buffer[64]<<2)+(in_buffer[64]<<4)+(in_buffer[64]<<5)+(in_buffer[64]<<8));
assign in_buffer_weight49=0+(0+(in_buffer[53]<<0)+(in_buffer[53]<<3)+(in_buffer[53]<<5)+(in_buffer[53]<<8))+(0+(in_buffer[54]<<1)+(in_buffer[54]<<2)+(in_buffer[54]<<8))+(0-(in_buffer[64]<<0)+(in_buffer[64]<<8))+(0+(in_buffer[65]<<2)+(in_buffer[65]<<4)+(in_buffer[65]<<5)+(in_buffer[65]<<8));
assign in_buffer_weight50=0+(0+(in_buffer[55]<<0)+(in_buffer[55]<<3)+(in_buffer[55]<<5)+(in_buffer[55]<<8))+(0+(in_buffer[56]<<1)+(in_buffer[56]<<2)+(in_buffer[56]<<8))+(0-(in_buffer[66]<<0)+(in_buffer[66]<<8))+(0+(in_buffer[67]<<2)+(in_buffer[67]<<4)+(in_buffer[67]<<5)+(in_buffer[67]<<8));
assign in_buffer_weight51=0+(0+(in_buffer[56]<<0)+(in_buffer[56]<<3)+(in_buffer[56]<<5)+(in_buffer[56]<<8))+(0+(in_buffer[57]<<1)+(in_buffer[57]<<2)+(in_buffer[57]<<8))+(0-(in_buffer[67]<<0)+(in_buffer[67]<<8))+(0+(in_buffer[68]<<2)+(in_buffer[68]<<4)+(in_buffer[68]<<5)+(in_buffer[68]<<8));
assign in_buffer_weight52=0+(0+(in_buffer[57]<<0)+(in_buffer[57]<<3)+(in_buffer[57]<<5)+(in_buffer[57]<<8))+(0+(in_buffer[58]<<1)+(in_buffer[58]<<2)+(in_buffer[58]<<8))+(0-(in_buffer[68]<<0)+(in_buffer[68]<<8))+(0+(in_buffer[69]<<2)+(in_buffer[69]<<4)+(in_buffer[69]<<5)+(in_buffer[69]<<8));
assign in_buffer_weight53=0+(0+(in_buffer[58]<<0)+(in_buffer[58]<<3)+(in_buffer[58]<<5)+(in_buffer[58]<<8))+(0+(in_buffer[59]<<1)+(in_buffer[59]<<2)+(in_buffer[59]<<8))+(0-(in_buffer[69]<<0)+(in_buffer[69]<<8))+(0+(in_buffer[70]<<2)+(in_buffer[70]<<4)+(in_buffer[70]<<5)+(in_buffer[70]<<8));
assign in_buffer_weight54=0+(0+(in_buffer[59]<<0)+(in_buffer[59]<<3)+(in_buffer[59]<<5)+(in_buffer[59]<<8))+(0+(in_buffer[60]<<1)+(in_buffer[60]<<2)+(in_buffer[60]<<8))+(0-(in_buffer[70]<<0)+(in_buffer[70]<<8))+(0+(in_buffer[71]<<2)+(in_buffer[71]<<4)+(in_buffer[71]<<5)+(in_buffer[71]<<8));
assign in_buffer_weight55=0+(0+(in_buffer[60]<<0)+(in_buffer[60]<<3)+(in_buffer[60]<<5)+(in_buffer[60]<<8))+(0+(in_buffer[61]<<1)+(in_buffer[61]<<2)+(in_buffer[61]<<8))+(0-(in_buffer[71]<<0)+(in_buffer[71]<<8))+(0+(in_buffer[72]<<2)+(in_buffer[72]<<4)+(in_buffer[72]<<5)+(in_buffer[72]<<8));
assign in_buffer_weight56=0+(0+(in_buffer[61]<<0)+(in_buffer[61]<<3)+(in_buffer[61]<<5)+(in_buffer[61]<<8))+(0+(in_buffer[62]<<1)+(in_buffer[62]<<2)+(in_buffer[62]<<8))+(0-(in_buffer[72]<<0)+(in_buffer[72]<<8))+(0+(in_buffer[73]<<2)+(in_buffer[73]<<4)+(in_buffer[73]<<5)+(in_buffer[73]<<8));
assign in_buffer_weight57=0+(0+(in_buffer[62]<<0)+(in_buffer[62]<<3)+(in_buffer[62]<<5)+(in_buffer[62]<<8))+(0+(in_buffer[63]<<1)+(in_buffer[63]<<2)+(in_buffer[63]<<8))+(0-(in_buffer[73]<<0)+(in_buffer[73]<<8))+(0+(in_buffer[74]<<2)+(in_buffer[74]<<4)+(in_buffer[74]<<5)+(in_buffer[74]<<8));
assign in_buffer_weight58=0+(0+(in_buffer[63]<<0)+(in_buffer[63]<<3)+(in_buffer[63]<<5)+(in_buffer[63]<<8))+(0+(in_buffer[64]<<1)+(in_buffer[64]<<2)+(in_buffer[64]<<8))+(0-(in_buffer[74]<<0)+(in_buffer[74]<<8))+(0+(in_buffer[75]<<2)+(in_buffer[75]<<4)+(in_buffer[75]<<5)+(in_buffer[75]<<8));
assign in_buffer_weight59=0+(0+(in_buffer[64]<<0)+(in_buffer[64]<<3)+(in_buffer[64]<<5)+(in_buffer[64]<<8))+(0+(in_buffer[65]<<1)+(in_buffer[65]<<2)+(in_buffer[65]<<8))+(0-(in_buffer[75]<<0)+(in_buffer[75]<<8))+(0+(in_buffer[76]<<2)+(in_buffer[76]<<4)+(in_buffer[76]<<5)+(in_buffer[76]<<8));
assign in_buffer_weight60=0+(0+(in_buffer[66]<<0)+(in_buffer[66]<<3)+(in_buffer[66]<<5)+(in_buffer[66]<<8))+(0+(in_buffer[67]<<1)+(in_buffer[67]<<2)+(in_buffer[67]<<8))+(0-(in_buffer[77]<<0)+(in_buffer[77]<<8))+(0+(in_buffer[78]<<2)+(in_buffer[78]<<4)+(in_buffer[78]<<5)+(in_buffer[78]<<8));
assign in_buffer_weight61=0+(0+(in_buffer[67]<<0)+(in_buffer[67]<<3)+(in_buffer[67]<<5)+(in_buffer[67]<<8))+(0+(in_buffer[68]<<1)+(in_buffer[68]<<2)+(in_buffer[68]<<8))+(0-(in_buffer[78]<<0)+(in_buffer[78]<<8))+(0+(in_buffer[79]<<2)+(in_buffer[79]<<4)+(in_buffer[79]<<5)+(in_buffer[79]<<8));
assign in_buffer_weight62=0+(0+(in_buffer[68]<<0)+(in_buffer[68]<<3)+(in_buffer[68]<<5)+(in_buffer[68]<<8))+(0+(in_buffer[69]<<1)+(in_buffer[69]<<2)+(in_buffer[69]<<8))+(0-(in_buffer[79]<<0)+(in_buffer[79]<<8))+(0+(in_buffer[80]<<2)+(in_buffer[80]<<4)+(in_buffer[80]<<5)+(in_buffer[80]<<8));
assign in_buffer_weight63=0+(0+(in_buffer[69]<<0)+(in_buffer[69]<<3)+(in_buffer[69]<<5)+(in_buffer[69]<<8))+(0+(in_buffer[70]<<1)+(in_buffer[70]<<2)+(in_buffer[70]<<8))+(0-(in_buffer[80]<<0)+(in_buffer[80]<<8))+(0+(in_buffer[81]<<2)+(in_buffer[81]<<4)+(in_buffer[81]<<5)+(in_buffer[81]<<8));
assign in_buffer_weight64=0+(0+(in_buffer[70]<<0)+(in_buffer[70]<<3)+(in_buffer[70]<<5)+(in_buffer[70]<<8))+(0+(in_buffer[71]<<1)+(in_buffer[71]<<2)+(in_buffer[71]<<8))+(0-(in_buffer[81]<<0)+(in_buffer[81]<<8))+(0+(in_buffer[82]<<2)+(in_buffer[82]<<4)+(in_buffer[82]<<5)+(in_buffer[82]<<8));
assign in_buffer_weight65=0+(0+(in_buffer[71]<<0)+(in_buffer[71]<<3)+(in_buffer[71]<<5)+(in_buffer[71]<<8))+(0+(in_buffer[72]<<1)+(in_buffer[72]<<2)+(in_buffer[72]<<8))+(0-(in_buffer[82]<<0)+(in_buffer[82]<<8))+(0+(in_buffer[83]<<2)+(in_buffer[83]<<4)+(in_buffer[83]<<5)+(in_buffer[83]<<8));
assign in_buffer_weight66=0+(0+(in_buffer[72]<<0)+(in_buffer[72]<<3)+(in_buffer[72]<<5)+(in_buffer[72]<<8))+(0+(in_buffer[73]<<1)+(in_buffer[73]<<2)+(in_buffer[73]<<8))+(0-(in_buffer[83]<<0)+(in_buffer[83]<<8))+(0+(in_buffer[84]<<2)+(in_buffer[84]<<4)+(in_buffer[84]<<5)+(in_buffer[84]<<8));
assign in_buffer_weight67=0+(0+(in_buffer[73]<<0)+(in_buffer[73]<<3)+(in_buffer[73]<<5)+(in_buffer[73]<<8))+(0+(in_buffer[74]<<1)+(in_buffer[74]<<2)+(in_buffer[74]<<8))+(0-(in_buffer[84]<<0)+(in_buffer[84]<<8))+(0+(in_buffer[85]<<2)+(in_buffer[85]<<4)+(in_buffer[85]<<5)+(in_buffer[85]<<8));
assign in_buffer_weight68=0+(0+(in_buffer[74]<<0)+(in_buffer[74]<<3)+(in_buffer[74]<<5)+(in_buffer[74]<<8))+(0+(in_buffer[75]<<1)+(in_buffer[75]<<2)+(in_buffer[75]<<8))+(0-(in_buffer[85]<<0)+(in_buffer[85]<<8))+(0+(in_buffer[86]<<2)+(in_buffer[86]<<4)+(in_buffer[86]<<5)+(in_buffer[86]<<8));
assign in_buffer_weight69=0+(0+(in_buffer[75]<<0)+(in_buffer[75]<<3)+(in_buffer[75]<<5)+(in_buffer[75]<<8))+(0+(in_buffer[76]<<1)+(in_buffer[76]<<2)+(in_buffer[76]<<8))+(0-(in_buffer[86]<<0)+(in_buffer[86]<<8))+(0+(in_buffer[87]<<2)+(in_buffer[87]<<4)+(in_buffer[87]<<5)+(in_buffer[87]<<8));
assign in_buffer_weight70=0+(0+(in_buffer[77]<<0)+(in_buffer[77]<<3)+(in_buffer[77]<<5)+(in_buffer[77]<<8))+(0+(in_buffer[78]<<1)+(in_buffer[78]<<2)+(in_buffer[78]<<8))+(0-(in_buffer[88]<<0)+(in_buffer[88]<<8))+(0+(in_buffer[89]<<2)+(in_buffer[89]<<4)+(in_buffer[89]<<5)+(in_buffer[89]<<8));
assign in_buffer_weight71=0+(0+(in_buffer[78]<<0)+(in_buffer[78]<<3)+(in_buffer[78]<<5)+(in_buffer[78]<<8))+(0+(in_buffer[79]<<1)+(in_buffer[79]<<2)+(in_buffer[79]<<8))+(0-(in_buffer[89]<<0)+(in_buffer[89]<<8))+(0+(in_buffer[90]<<2)+(in_buffer[90]<<4)+(in_buffer[90]<<5)+(in_buffer[90]<<8));
assign in_buffer_weight72=0+(0+(in_buffer[79]<<0)+(in_buffer[79]<<3)+(in_buffer[79]<<5)+(in_buffer[79]<<8))+(0+(in_buffer[80]<<1)+(in_buffer[80]<<2)+(in_buffer[80]<<8))+(0-(in_buffer[90]<<0)+(in_buffer[90]<<8))+(0+(in_buffer[91]<<2)+(in_buffer[91]<<4)+(in_buffer[91]<<5)+(in_buffer[91]<<8));
assign in_buffer_weight73=0+(0+(in_buffer[80]<<0)+(in_buffer[80]<<3)+(in_buffer[80]<<5)+(in_buffer[80]<<8))+(0+(in_buffer[81]<<1)+(in_buffer[81]<<2)+(in_buffer[81]<<8))+(0-(in_buffer[91]<<0)+(in_buffer[91]<<8))+(0+(in_buffer[92]<<2)+(in_buffer[92]<<4)+(in_buffer[92]<<5)+(in_buffer[92]<<8));
assign in_buffer_weight74=0+(0+(in_buffer[81]<<0)+(in_buffer[81]<<3)+(in_buffer[81]<<5)+(in_buffer[81]<<8))+(0+(in_buffer[82]<<1)+(in_buffer[82]<<2)+(in_buffer[82]<<8))+(0-(in_buffer[92]<<0)+(in_buffer[92]<<8))+(0+(in_buffer[93]<<2)+(in_buffer[93]<<4)+(in_buffer[93]<<5)+(in_buffer[93]<<8));
assign in_buffer_weight75=0+(0+(in_buffer[82]<<0)+(in_buffer[82]<<3)+(in_buffer[82]<<5)+(in_buffer[82]<<8))+(0+(in_buffer[83]<<1)+(in_buffer[83]<<2)+(in_buffer[83]<<8))+(0-(in_buffer[93]<<0)+(in_buffer[93]<<8))+(0+(in_buffer[94]<<2)+(in_buffer[94]<<4)+(in_buffer[94]<<5)+(in_buffer[94]<<8));
assign in_buffer_weight76=0+(0+(in_buffer[83]<<0)+(in_buffer[83]<<3)+(in_buffer[83]<<5)+(in_buffer[83]<<8))+(0+(in_buffer[84]<<1)+(in_buffer[84]<<2)+(in_buffer[84]<<8))+(0-(in_buffer[94]<<0)+(in_buffer[94]<<8))+(0+(in_buffer[95]<<2)+(in_buffer[95]<<4)+(in_buffer[95]<<5)+(in_buffer[95]<<8));
assign in_buffer_weight77=0+(0+(in_buffer[84]<<0)+(in_buffer[84]<<3)+(in_buffer[84]<<5)+(in_buffer[84]<<8))+(0+(in_buffer[85]<<1)+(in_buffer[85]<<2)+(in_buffer[85]<<8))+(0-(in_buffer[95]<<0)+(in_buffer[95]<<8))+(0+(in_buffer[96]<<2)+(in_buffer[96]<<4)+(in_buffer[96]<<5)+(in_buffer[96]<<8));
assign in_buffer_weight78=0+(0+(in_buffer[85]<<0)+(in_buffer[85]<<3)+(in_buffer[85]<<5)+(in_buffer[85]<<8))+(0+(in_buffer[86]<<1)+(in_buffer[86]<<2)+(in_buffer[86]<<8))+(0-(in_buffer[96]<<0)+(in_buffer[96]<<8))+(0+(in_buffer[97]<<2)+(in_buffer[97]<<4)+(in_buffer[97]<<5)+(in_buffer[97]<<8));
assign in_buffer_weight79=0+(0+(in_buffer[86]<<0)+(in_buffer[86]<<3)+(in_buffer[86]<<5)+(in_buffer[86]<<8))+(0+(in_buffer[87]<<1)+(in_buffer[87]<<2)+(in_buffer[87]<<8))+(0-(in_buffer[97]<<0)+(in_buffer[97]<<8))+(0+(in_buffer[98]<<2)+(in_buffer[98]<<4)+(in_buffer[98]<<5)+(in_buffer[98]<<8));
assign in_buffer_weight80=0+(0+(in_buffer[88]<<0)+(in_buffer[88]<<3)+(in_buffer[88]<<5)+(in_buffer[88]<<8))+(0+(in_buffer[89]<<1)+(in_buffer[89]<<2)+(in_buffer[89]<<8))+(0-(in_buffer[99]<<0)+(in_buffer[99]<<8))+(0+(in_buffer[100]<<2)+(in_buffer[100]<<4)+(in_buffer[100]<<5)+(in_buffer[100]<<8));
assign in_buffer_weight81=0+(0+(in_buffer[89]<<0)+(in_buffer[89]<<3)+(in_buffer[89]<<5)+(in_buffer[89]<<8))+(0+(in_buffer[90]<<1)+(in_buffer[90]<<2)+(in_buffer[90]<<8))+(0-(in_buffer[100]<<0)+(in_buffer[100]<<8))+(0+(in_buffer[101]<<2)+(in_buffer[101]<<4)+(in_buffer[101]<<5)+(in_buffer[101]<<8));
assign in_buffer_weight82=0+(0+(in_buffer[90]<<0)+(in_buffer[90]<<3)+(in_buffer[90]<<5)+(in_buffer[90]<<8))+(0+(in_buffer[91]<<1)+(in_buffer[91]<<2)+(in_buffer[91]<<8))+(0-(in_buffer[101]<<0)+(in_buffer[101]<<8))+(0+(in_buffer[102]<<2)+(in_buffer[102]<<4)+(in_buffer[102]<<5)+(in_buffer[102]<<8));
assign in_buffer_weight83=0+(0+(in_buffer[91]<<0)+(in_buffer[91]<<3)+(in_buffer[91]<<5)+(in_buffer[91]<<8))+(0+(in_buffer[92]<<1)+(in_buffer[92]<<2)+(in_buffer[92]<<8))+(0-(in_buffer[102]<<0)+(in_buffer[102]<<8))+(0+(in_buffer[103]<<2)+(in_buffer[103]<<4)+(in_buffer[103]<<5)+(in_buffer[103]<<8));
assign in_buffer_weight84=0+(0+(in_buffer[92]<<0)+(in_buffer[92]<<3)+(in_buffer[92]<<5)+(in_buffer[92]<<8))+(0+(in_buffer[93]<<1)+(in_buffer[93]<<2)+(in_buffer[93]<<8))+(0-(in_buffer[103]<<0)+(in_buffer[103]<<8))+(0+(in_buffer[104]<<2)+(in_buffer[104]<<4)+(in_buffer[104]<<5)+(in_buffer[104]<<8));
assign in_buffer_weight85=0+(0+(in_buffer[93]<<0)+(in_buffer[93]<<3)+(in_buffer[93]<<5)+(in_buffer[93]<<8))+(0+(in_buffer[94]<<1)+(in_buffer[94]<<2)+(in_buffer[94]<<8))+(0-(in_buffer[104]<<0)+(in_buffer[104]<<8))+(0+(in_buffer[105]<<2)+(in_buffer[105]<<4)+(in_buffer[105]<<5)+(in_buffer[105]<<8));
assign in_buffer_weight86=0+(0+(in_buffer[94]<<0)+(in_buffer[94]<<3)+(in_buffer[94]<<5)+(in_buffer[94]<<8))+(0+(in_buffer[95]<<1)+(in_buffer[95]<<2)+(in_buffer[95]<<8))+(0-(in_buffer[105]<<0)+(in_buffer[105]<<8))+(0+(in_buffer[106]<<2)+(in_buffer[106]<<4)+(in_buffer[106]<<5)+(in_buffer[106]<<8));
assign in_buffer_weight87=0+(0+(in_buffer[95]<<0)+(in_buffer[95]<<3)+(in_buffer[95]<<5)+(in_buffer[95]<<8))+(0+(in_buffer[96]<<1)+(in_buffer[96]<<2)+(in_buffer[96]<<8))+(0-(in_buffer[106]<<0)+(in_buffer[106]<<8))+(0+(in_buffer[107]<<2)+(in_buffer[107]<<4)+(in_buffer[107]<<5)+(in_buffer[107]<<8));
assign in_buffer_weight88=0+(0+(in_buffer[96]<<0)+(in_buffer[96]<<3)+(in_buffer[96]<<5)+(in_buffer[96]<<8))+(0+(in_buffer[97]<<1)+(in_buffer[97]<<2)+(in_buffer[97]<<8))+(0-(in_buffer[107]<<0)+(in_buffer[107]<<8))+(0+(in_buffer[108]<<2)+(in_buffer[108]<<4)+(in_buffer[108]<<5)+(in_buffer[108]<<8));
assign in_buffer_weight89=0+(0+(in_buffer[97]<<0)+(in_buffer[97]<<3)+(in_buffer[97]<<5)+(in_buffer[97]<<8))+(0+(in_buffer[98]<<1)+(in_buffer[98]<<2)+(in_buffer[98]<<8))+(0-(in_buffer[108]<<0)+(in_buffer[108]<<8))+(0+(in_buffer[109]<<2)+(in_buffer[109]<<4)+(in_buffer[109]<<5)+(in_buffer[109]<<8));
assign in_buffer_weight90=0+(0+(in_buffer[99]<<0)+(in_buffer[99]<<3)+(in_buffer[99]<<5)+(in_buffer[99]<<8))+(0+(in_buffer[100]<<1)+(in_buffer[100]<<2)+(in_buffer[100]<<8))+(0-(in_buffer[110]<<0)+(in_buffer[110]<<8))+(0+(in_buffer[111]<<2)+(in_buffer[111]<<4)+(in_buffer[111]<<5)+(in_buffer[111]<<8));
assign in_buffer_weight91=0+(0+(in_buffer[100]<<0)+(in_buffer[100]<<3)+(in_buffer[100]<<5)+(in_buffer[100]<<8))+(0+(in_buffer[101]<<1)+(in_buffer[101]<<2)+(in_buffer[101]<<8))+(0-(in_buffer[111]<<0)+(in_buffer[111]<<8))+(0+(in_buffer[112]<<2)+(in_buffer[112]<<4)+(in_buffer[112]<<5)+(in_buffer[112]<<8));
assign in_buffer_weight92=0+(0+(in_buffer[101]<<0)+(in_buffer[101]<<3)+(in_buffer[101]<<5)+(in_buffer[101]<<8))+(0+(in_buffer[102]<<1)+(in_buffer[102]<<2)+(in_buffer[102]<<8))+(0-(in_buffer[112]<<0)+(in_buffer[112]<<8))+(0+(in_buffer[113]<<2)+(in_buffer[113]<<4)+(in_buffer[113]<<5)+(in_buffer[113]<<8));
assign in_buffer_weight93=0+(0+(in_buffer[102]<<0)+(in_buffer[102]<<3)+(in_buffer[102]<<5)+(in_buffer[102]<<8))+(0+(in_buffer[103]<<1)+(in_buffer[103]<<2)+(in_buffer[103]<<8))+(0-(in_buffer[113]<<0)+(in_buffer[113]<<8))+(0+(in_buffer[114]<<2)+(in_buffer[114]<<4)+(in_buffer[114]<<5)+(in_buffer[114]<<8));
assign in_buffer_weight94=0+(0+(in_buffer[103]<<0)+(in_buffer[103]<<3)+(in_buffer[103]<<5)+(in_buffer[103]<<8))+(0+(in_buffer[104]<<1)+(in_buffer[104]<<2)+(in_buffer[104]<<8))+(0-(in_buffer[114]<<0)+(in_buffer[114]<<8))+(0+(in_buffer[115]<<2)+(in_buffer[115]<<4)+(in_buffer[115]<<5)+(in_buffer[115]<<8));
assign in_buffer_weight95=0+(0+(in_buffer[104]<<0)+(in_buffer[104]<<3)+(in_buffer[104]<<5)+(in_buffer[104]<<8))+(0+(in_buffer[105]<<1)+(in_buffer[105]<<2)+(in_buffer[105]<<8))+(0-(in_buffer[115]<<0)+(in_buffer[115]<<8))+(0+(in_buffer[116]<<2)+(in_buffer[116]<<4)+(in_buffer[116]<<5)+(in_buffer[116]<<8));
assign in_buffer_weight96=0+(0+(in_buffer[105]<<0)+(in_buffer[105]<<3)+(in_buffer[105]<<5)+(in_buffer[105]<<8))+(0+(in_buffer[106]<<1)+(in_buffer[106]<<2)+(in_buffer[106]<<8))+(0-(in_buffer[116]<<0)+(in_buffer[116]<<8))+(0+(in_buffer[117]<<2)+(in_buffer[117]<<4)+(in_buffer[117]<<5)+(in_buffer[117]<<8));
assign in_buffer_weight97=0+(0+(in_buffer[106]<<0)+(in_buffer[106]<<3)+(in_buffer[106]<<5)+(in_buffer[106]<<8))+(0+(in_buffer[107]<<1)+(in_buffer[107]<<2)+(in_buffer[107]<<8))+(0-(in_buffer[117]<<0)+(in_buffer[117]<<8))+(0+(in_buffer[118]<<2)+(in_buffer[118]<<4)+(in_buffer[118]<<5)+(in_buffer[118]<<8));
assign in_buffer_weight98=0+(0+(in_buffer[107]<<0)+(in_buffer[107]<<3)+(in_buffer[107]<<5)+(in_buffer[107]<<8))+(0+(in_buffer[108]<<1)+(in_buffer[108]<<2)+(in_buffer[108]<<8))+(0-(in_buffer[118]<<0)+(in_buffer[118]<<8))+(0+(in_buffer[119]<<2)+(in_buffer[119]<<4)+(in_buffer[119]<<5)+(in_buffer[119]<<8));
assign in_buffer_weight99=0+(0+(in_buffer[108]<<0)+(in_buffer[108]<<3)+(in_buffer[108]<<5)+(in_buffer[108]<<8))+(0+(in_buffer[109]<<1)+(in_buffer[109]<<2)+(in_buffer[109]<<8))+(0-(in_buffer[119]<<0)+(in_buffer[119]<<8))+(0+(in_buffer[120]<<2)+(in_buffer[120]<<4)+(in_buffer[120]<<5)+(in_buffer[120]<<8));
wire signed    [DATA_WIDTH-1:0]   weight_bias0;
assign weight_bias0= in_buffer_weight0+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias1;
assign weight_bias1= in_buffer_weight1+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias2;
assign weight_bias2= in_buffer_weight2+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias3;
assign weight_bias3= in_buffer_weight3+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias4;
assign weight_bias4= in_buffer_weight4+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias5;
assign weight_bias5= in_buffer_weight5+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias6;
assign weight_bias6= in_buffer_weight6+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias7;
assign weight_bias7= in_buffer_weight7+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias8;
assign weight_bias8= in_buffer_weight8+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias9= in_buffer_weight9+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias10;
assign weight_bias10= in_buffer_weight10+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias11;
assign weight_bias11= in_buffer_weight11+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias12;
assign weight_bias12= in_buffer_weight12+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias13;
assign weight_bias13= in_buffer_weight13+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias14;
assign weight_bias14= in_buffer_weight14+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias15;
assign weight_bias15= in_buffer_weight15+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias16;
assign weight_bias16= in_buffer_weight16+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias17;
assign weight_bias17= in_buffer_weight17+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias18;
assign weight_bias18= in_buffer_weight18+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias19;
assign weight_bias19= in_buffer_weight19+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias20;
assign weight_bias20= in_buffer_weight20+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias21;
assign weight_bias21= in_buffer_weight21+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias22;
assign weight_bias22= in_buffer_weight22+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias23;
assign weight_bias23= in_buffer_weight23+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias24;
assign weight_bias24= in_buffer_weight24+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias25;
assign weight_bias25= in_buffer_weight25+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias26;
assign weight_bias26= in_buffer_weight26+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias27;
assign weight_bias27= in_buffer_weight27+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias28;
assign weight_bias28= in_buffer_weight28+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias29;
assign weight_bias29= in_buffer_weight29+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias30;
assign weight_bias30= in_buffer_weight30+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias31;
assign weight_bias31= in_buffer_weight31+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias32;
assign weight_bias32= in_buffer_weight32+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias33;
assign weight_bias33= in_buffer_weight33+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias34;
assign weight_bias34= in_buffer_weight34+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias35;
assign weight_bias35= in_buffer_weight35+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias36;
assign weight_bias36= in_buffer_weight36+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias37;
assign weight_bias37= in_buffer_weight37+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias38;
assign weight_bias38= in_buffer_weight38+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias39;
assign weight_bias39= in_buffer_weight39+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias40;
assign weight_bias40= in_buffer_weight40+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias41;
assign weight_bias41= in_buffer_weight41+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias42;
assign weight_bias42= in_buffer_weight42+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias43;
assign weight_bias43= in_buffer_weight43+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias44;
assign weight_bias44= in_buffer_weight44+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias45;
assign weight_bias45= in_buffer_weight45+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias46;
assign weight_bias46= in_buffer_weight46+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias47;
assign weight_bias47= in_buffer_weight47+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias48;
assign weight_bias48= in_buffer_weight48+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias49;
assign weight_bias49= in_buffer_weight49+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias50;
assign weight_bias50= in_buffer_weight50+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias51;
assign weight_bias51= in_buffer_weight51+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias52;
assign weight_bias52= in_buffer_weight52+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias53;
assign weight_bias53= in_buffer_weight53+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias54;
assign weight_bias54= in_buffer_weight54+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias55;
assign weight_bias55= in_buffer_weight55+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias56;
assign weight_bias56= in_buffer_weight56+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias57;
assign weight_bias57= in_buffer_weight57+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias58;
assign weight_bias58= in_buffer_weight58+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias59;
assign weight_bias59= in_buffer_weight59+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias60;
assign weight_bias60= in_buffer_weight60+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias61;
assign weight_bias61= in_buffer_weight61+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias62;
assign weight_bias62= in_buffer_weight62+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias63;
assign weight_bias63= in_buffer_weight63+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias64;
assign weight_bias64= in_buffer_weight64+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias65;
assign weight_bias65= in_buffer_weight65+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias66;
assign weight_bias66= in_buffer_weight66+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias67;
assign weight_bias67= in_buffer_weight67+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias68;
assign weight_bias68= in_buffer_weight68+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias69;
assign weight_bias69= in_buffer_weight69+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias70;
assign weight_bias70= in_buffer_weight70+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias71;
assign weight_bias71= in_buffer_weight71+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias72;
assign weight_bias72= in_buffer_weight72+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias73;
assign weight_bias73= in_buffer_weight73+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias74;
assign weight_bias74= in_buffer_weight74+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias75;
assign weight_bias75= in_buffer_weight75+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias76;
assign weight_bias76= in_buffer_weight76+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias77;
assign weight_bias77= in_buffer_weight77+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias78;
assign weight_bias78= in_buffer_weight78+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias79;
assign weight_bias79= in_buffer_weight79+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias80;
assign weight_bias80= in_buffer_weight80+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias81;
assign weight_bias81= in_buffer_weight81+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias82;
assign weight_bias82= in_buffer_weight82+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias83;
assign weight_bias83= in_buffer_weight83+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias84;
assign weight_bias84= in_buffer_weight84+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias85;
assign weight_bias85= in_buffer_weight85+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias86;
assign weight_bias86= in_buffer_weight86+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias87;
assign weight_bias87= in_buffer_weight87+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias88;
assign weight_bias88= in_buffer_weight88+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias89;
assign weight_bias89= in_buffer_weight89+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias90;
assign weight_bias90= in_buffer_weight90+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias91;
assign weight_bias91= in_buffer_weight91+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias92;
assign weight_bias92= in_buffer_weight92+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias93;
assign weight_bias93= in_buffer_weight93+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias94;
assign weight_bias94= in_buffer_weight94+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias95;
assign weight_bias95= in_buffer_weight95+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias96;
assign weight_bias96= in_buffer_weight96+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias97;
assign weight_bias97= in_buffer_weight97+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias98;
assign weight_bias98= in_buffer_weight98+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias99;
assign weight_bias99= in_buffer_weight99+1;
wire signed    [DATA_WIDTH-1:0]   bias_relu0;
wire signed    [DATA_WIDTH-1:0]   bias_relu1;
wire signed    [DATA_WIDTH-1:0]   bias_relu2;
wire signed    [DATA_WIDTH-1:0]   bias_relu3;
wire signed    [DATA_WIDTH-1:0]   bias_relu4;
wire signed    [DATA_WIDTH-1:0]   bias_relu5;
wire signed    [DATA_WIDTH-1:0]   bias_relu6;
wire signed    [DATA_WIDTH-1:0]   bias_relu7;
wire signed    [DATA_WIDTH-1:0]   bias_relu8;
wire signed    [DATA_WIDTH-1:0]   bias_relu9;
wire signed    [DATA_WIDTH-1:0]   bias_relu10;
wire signed    [DATA_WIDTH-1:0]   bias_relu11;
wire signed    [DATA_WIDTH-1:0]   bias_relu12;
wire signed    [DATA_WIDTH-1:0]   bias_relu13;
wire signed    [DATA_WIDTH-1:0]   bias_relu14;
wire signed    [DATA_WIDTH-1:0]   bias_relu15;
wire signed    [DATA_WIDTH-1:0]   bias_relu16;
wire signed    [DATA_WIDTH-1:0]   bias_relu17;
wire signed    [DATA_WIDTH-1:0]   bias_relu18;
wire signed    [DATA_WIDTH-1:0]   bias_relu19;
wire signed    [DATA_WIDTH-1:0]   bias_relu20;
wire signed    [DATA_WIDTH-1:0]   bias_relu21;
wire signed    [DATA_WIDTH-1:0]   bias_relu22;
wire signed    [DATA_WIDTH-1:0]   bias_relu23;
wire signed    [DATA_WIDTH-1:0]   bias_relu24;
wire signed    [DATA_WIDTH-1:0]   bias_relu25;
wire signed    [DATA_WIDTH-1:0]   bias_relu26;
wire signed    [DATA_WIDTH-1:0]   bias_relu27;
wire signed    [DATA_WIDTH-1:0]   bias_relu28;
wire signed    [DATA_WIDTH-1:0]   bias_relu29;
wire signed    [DATA_WIDTH-1:0]   bias_relu30;
wire signed    [DATA_WIDTH-1:0]   bias_relu31;
wire signed    [DATA_WIDTH-1:0]   bias_relu32;
wire signed    [DATA_WIDTH-1:0]   bias_relu33;
wire signed    [DATA_WIDTH-1:0]   bias_relu34;
wire signed    [DATA_WIDTH-1:0]   bias_relu35;
wire signed    [DATA_WIDTH-1:0]   bias_relu36;
wire signed    [DATA_WIDTH-1:0]   bias_relu37;
wire signed    [DATA_WIDTH-1:0]   bias_relu38;
wire signed    [DATA_WIDTH-1:0]   bias_relu39;
wire signed    [DATA_WIDTH-1:0]   bias_relu40;
wire signed    [DATA_WIDTH-1:0]   bias_relu41;
wire signed    [DATA_WIDTH-1:0]   bias_relu42;
wire signed    [DATA_WIDTH-1:0]   bias_relu43;
wire signed    [DATA_WIDTH-1:0]   bias_relu44;
wire signed    [DATA_WIDTH-1:0]   bias_relu45;
wire signed    [DATA_WIDTH-1:0]   bias_relu46;
wire signed    [DATA_WIDTH-1:0]   bias_relu47;
wire signed    [DATA_WIDTH-1:0]   bias_relu48;
wire signed    [DATA_WIDTH-1:0]   bias_relu49;
wire signed    [DATA_WIDTH-1:0]   bias_relu50;
wire signed    [DATA_WIDTH-1:0]   bias_relu51;
wire signed    [DATA_WIDTH-1:0]   bias_relu52;
wire signed    [DATA_WIDTH-1:0]   bias_relu53;
wire signed    [DATA_WIDTH-1:0]   bias_relu54;
wire signed    [DATA_WIDTH-1:0]   bias_relu55;
wire signed    [DATA_WIDTH-1:0]   bias_relu56;
wire signed    [DATA_WIDTH-1:0]   bias_relu57;
wire signed    [DATA_WIDTH-1:0]   bias_relu58;
wire signed    [DATA_WIDTH-1:0]   bias_relu59;
wire signed    [DATA_WIDTH-1:0]   bias_relu60;
wire signed    [DATA_WIDTH-1:0]   bias_relu61;
wire signed    [DATA_WIDTH-1:0]   bias_relu62;
wire signed    [DATA_WIDTH-1:0]   bias_relu63;
wire signed    [DATA_WIDTH-1:0]   bias_relu64;
wire signed    [DATA_WIDTH-1:0]   bias_relu65;
wire signed    [DATA_WIDTH-1:0]   bias_relu66;
wire signed    [DATA_WIDTH-1:0]   bias_relu67;
wire signed    [DATA_WIDTH-1:0]   bias_relu68;
wire signed    [DATA_WIDTH-1:0]   bias_relu69;
wire signed    [DATA_WIDTH-1:0]   bias_relu70;
wire signed    [DATA_WIDTH-1:0]   bias_relu71;
wire signed    [DATA_WIDTH-1:0]   bias_relu72;
wire signed    [DATA_WIDTH-1:0]   bias_relu73;
wire signed    [DATA_WIDTH-1:0]   bias_relu74;
wire signed    [DATA_WIDTH-1:0]   bias_relu75;
wire signed    [DATA_WIDTH-1:0]   bias_relu76;
wire signed    [DATA_WIDTH-1:0]   bias_relu77;
wire signed    [DATA_WIDTH-1:0]   bias_relu78;
wire signed    [DATA_WIDTH-1:0]   bias_relu79;
wire signed    [DATA_WIDTH-1:0]   bias_relu80;
wire signed    [DATA_WIDTH-1:0]   bias_relu81;
wire signed    [DATA_WIDTH-1:0]   bias_relu82;
wire signed    [DATA_WIDTH-1:0]   bias_relu83;
wire signed    [DATA_WIDTH-1:0]   bias_relu84;
wire signed    [DATA_WIDTH-1:0]   bias_relu85;
wire signed    [DATA_WIDTH-1:0]   bias_relu86;
wire signed    [DATA_WIDTH-1:0]   bias_relu87;
wire signed    [DATA_WIDTH-1:0]   bias_relu88;
wire signed    [DATA_WIDTH-1:0]   bias_relu89;
wire signed    [DATA_WIDTH-1:0]   bias_relu90;
wire signed    [DATA_WIDTH-1:0]   bias_relu91;
wire signed    [DATA_WIDTH-1:0]   bias_relu92;
wire signed    [DATA_WIDTH-1:0]   bias_relu93;
wire signed    [DATA_WIDTH-1:0]   bias_relu94;
wire signed    [DATA_WIDTH-1:0]   bias_relu95;
wire signed    [DATA_WIDTH-1:0]   bias_relu96;
wire signed    [DATA_WIDTH-1:0]   bias_relu97;
wire signed    [DATA_WIDTH-1:0]   bias_relu98;
wire signed    [DATA_WIDTH-1:0]   bias_relu99;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign bias_relu32=(weight_bias32[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias32;
assign bias_relu33=(weight_bias33[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias33;
assign bias_relu34=(weight_bias34[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias34;
assign bias_relu35=(weight_bias35[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias35;
assign bias_relu36=(weight_bias36[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias36;
assign bias_relu37=(weight_bias37[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias37;
assign bias_relu38=(weight_bias38[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias38;
assign bias_relu39=(weight_bias39[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias39;
assign bias_relu40=(weight_bias40[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias40;
assign bias_relu41=(weight_bias41[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias41;
assign bias_relu42=(weight_bias42[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias42;
assign bias_relu43=(weight_bias43[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias43;
assign bias_relu44=(weight_bias44[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias44;
assign bias_relu45=(weight_bias45[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias45;
assign bias_relu46=(weight_bias46[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias46;
assign bias_relu47=(weight_bias47[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias47;
assign bias_relu48=(weight_bias48[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias48;
assign bias_relu49=(weight_bias49[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias49;
assign bias_relu50=(weight_bias50[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias50;
assign bias_relu51=(weight_bias51[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias51;
assign bias_relu52=(weight_bias52[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias52;
assign bias_relu53=(weight_bias53[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias53;
assign bias_relu54=(weight_bias54[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias54;
assign bias_relu55=(weight_bias55[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias55;
assign bias_relu56=(weight_bias56[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias56;
assign bias_relu57=(weight_bias57[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias57;
assign bias_relu58=(weight_bias58[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias58;
assign bias_relu59=(weight_bias59[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias59;
assign bias_relu60=(weight_bias60[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias60;
assign bias_relu61=(weight_bias61[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias61;
assign bias_relu62=(weight_bias62[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias62;
assign bias_relu63=(weight_bias63[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias63;
assign bias_relu64=(weight_bias64[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias64;
assign bias_relu65=(weight_bias65[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias65;
assign bias_relu66=(weight_bias66[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias66;
assign bias_relu67=(weight_bias67[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias67;
assign bias_relu68=(weight_bias68[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias68;
assign bias_relu69=(weight_bias69[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias69;
assign bias_relu70=(weight_bias70[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias70;
assign bias_relu71=(weight_bias71[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias71;
assign bias_relu72=(weight_bias72[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias72;
assign bias_relu73=(weight_bias73[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias73;
assign bias_relu74=(weight_bias74[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias74;
assign bias_relu75=(weight_bias75[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias75;
assign bias_relu76=(weight_bias76[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias76;
assign bias_relu77=(weight_bias77[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias77;
assign bias_relu78=(weight_bias78[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias78;
assign bias_relu79=(weight_bias79[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias79;
assign bias_relu80=(weight_bias80[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias80;
assign bias_relu81=(weight_bias81[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias81;
assign bias_relu82=(weight_bias82[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias82;
assign bias_relu83=(weight_bias83[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias83;
assign bias_relu84=(weight_bias84[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias84;
assign bias_relu85=(weight_bias85[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias85;
assign bias_relu86=(weight_bias86[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias86;
assign bias_relu87=(weight_bias87[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias87;
assign bias_relu88=(weight_bias88[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias88;
assign bias_relu89=(weight_bias89[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias89;
assign bias_relu90=(weight_bias90[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias90;
assign bias_relu91=(weight_bias91[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias91;
assign bias_relu92=(weight_bias92[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias92;
assign bias_relu93=(weight_bias93[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias93;
assign bias_relu94=(weight_bias94[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias94;
assign bias_relu95=(weight_bias95[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias95;
assign bias_relu96=(weight_bias96[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias96;
assign bias_relu97=(weight_bias97[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias97;
assign bias_relu98=(weight_bias98[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias98;
assign bias_relu99=(weight_bias99[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias99;
assign layer_out={
bias_relu99,bias_relu98,bias_relu97,bias_relu96,bias_relu95,bias_relu94,bias_relu93,bias_relu92,bias_relu91,bias_relu90,bias_relu89,bias_relu88,bias_relu87,bias_relu86,bias_relu85,bias_relu84,bias_relu83,bias_relu82,bias_relu81,bias_relu80,bias_relu79,bias_relu78,bias_relu77,bias_relu76,bias_relu75,bias_relu74,bias_relu73,bias_relu72,bias_relu71,bias_relu70,bias_relu69,bias_relu68,bias_relu67,bias_relu66,bias_relu65,bias_relu64,bias_relu63,bias_relu62,bias_relu61,bias_relu60,bias_relu59,bias_relu58,bias_relu57,bias_relu56,bias_relu55,bias_relu54,bias_relu53,bias_relu52,bias_relu51,bias_relu50,bias_relu49,bias_relu48,bias_relu47,bias_relu46,bias_relu45,bias_relu44,bias_relu43,bias_relu42,bias_relu41,bias_relu40,bias_relu39,bias_relu38,bias_relu37,bias_relu36,bias_relu35,bias_relu34,bias_relu33,bias_relu32,bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule