module layer2_tcb_121x64x10
(
    input clk,
    input rst,
   input valid,
   output  reg ready,
    input [25*64-1:0]  layer_in,
    output [42*10-1:0]   layer_out
);
parameter DATA_WIDTH   =   42;
reg [DATA_WIDTH-1:0]    layer_in_buffer    [0:64-1];
integer i;
always@(posedge clk )
    begin
        if(rst)
            begin
                for(i=0;i<64;i=i+1)
                    begin
                        layer_in_buffer[i]<=0;
                    end
            end
        else
        begin
       layer_in_buffer[0]<=layer_in[24:0];
       layer_in_buffer[1]<=layer_in[49:25];
       layer_in_buffer[2]<=layer_in[74:50];
       layer_in_buffer[3]<=layer_in[99:75];
       layer_in_buffer[4]<=layer_in[124:100];
       layer_in_buffer[5]<=layer_in[149:125];
       layer_in_buffer[6]<=layer_in[174:150];
       layer_in_buffer[7]<=layer_in[199:175];
       layer_in_buffer[8]<=layer_in[224:200];
       layer_in_buffer[9]<=layer_in[249:225];
       layer_in_buffer[10]<=layer_in[274:250];
       layer_in_buffer[11]<=layer_in[299:275];
       layer_in_buffer[12]<=layer_in[324:300];
       layer_in_buffer[13]<=layer_in[349:325];
       layer_in_buffer[14]<=layer_in[374:350];
       layer_in_buffer[15]<=layer_in[399:375];
       layer_in_buffer[16]<=layer_in[424:400];
       layer_in_buffer[17]<=layer_in[449:425];
       layer_in_buffer[18]<=layer_in[474:450];
       layer_in_buffer[19]<=layer_in[499:475];
       layer_in_buffer[20]<=layer_in[524:500];
       layer_in_buffer[21]<=layer_in[549:525];
       layer_in_buffer[22]<=layer_in[574:550];
       layer_in_buffer[23]<=layer_in[599:575];
       layer_in_buffer[24]<=layer_in[624:600];
       layer_in_buffer[25]<=layer_in[649:625];
       layer_in_buffer[26]<=layer_in[674:650];
       layer_in_buffer[27]<=layer_in[699:675];
       layer_in_buffer[28]<=layer_in[724:700];
       layer_in_buffer[29]<=layer_in[749:725];
       layer_in_buffer[30]<=layer_in[774:750];
       layer_in_buffer[31]<=layer_in[799:775];
       layer_in_buffer[32]<=layer_in[824:800];
       layer_in_buffer[33]<=layer_in[849:825];
       layer_in_buffer[34]<=layer_in[874:850];
       layer_in_buffer[35]<=layer_in[899:875];
       layer_in_buffer[36]<=layer_in[924:900];
       layer_in_buffer[37]<=layer_in[949:925];
       layer_in_buffer[38]<=layer_in[974:950];
       layer_in_buffer[39]<=layer_in[999:975];
       layer_in_buffer[40]<=layer_in[1024:1000];
       layer_in_buffer[41]<=layer_in[1049:1025];
       layer_in_buffer[42]<=layer_in[1074:1050];
       layer_in_buffer[43]<=layer_in[1099:1075];
       layer_in_buffer[44]<=layer_in[1124:1100];
       layer_in_buffer[45]<=layer_in[1149:1125];
       layer_in_buffer[46]<=layer_in[1174:1150];
       layer_in_buffer[47]<=layer_in[1199:1175];
       layer_in_buffer[48]<=layer_in[1224:1200];
       layer_in_buffer[49]<=layer_in[1249:1225];
       layer_in_buffer[50]<=layer_in[1274:1250];
       layer_in_buffer[51]<=layer_in[1299:1275];
       layer_in_buffer[52]<=layer_in[1324:1300];
       layer_in_buffer[53]<=layer_in[1349:1325];
       layer_in_buffer[54]<=layer_in[1374:1350];
       layer_in_buffer[55]<=layer_in[1399:1375];
       layer_in_buffer[56]<=layer_in[1424:1400];
       layer_in_buffer[57]<=layer_in[1449:1425];
       layer_in_buffer[58]<=layer_in[1474:1450];
       layer_in_buffer[59]<=layer_in[1499:1475];
       layer_in_buffer[60]<=layer_in[1524:1500];
       layer_in_buffer[61]<=layer_in[1549:1525];
       layer_in_buffer[62]<=layer_in[1574:1550];
       layer_in_buffer[63]<=layer_in[1599:1575];
        end
   end

wire [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0-(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)-(layer_in_buffer[0]<<5)+(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<10))-(0+(layer_in_buffer[1]<<0)+(layer_in_buffer[1]<<1)-(layer_in_buffer[1]<<4)-(layer_in_buffer[1]<<6)-(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<10)+(layer_in_buffer[1]<<11))-(0+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<7)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<12))+(0+(layer_in_buffer[3]<<1)+(layer_in_buffer[3]<<2)-(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<11))+(0+(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<11)+(layer_in_buffer[4]<<13))-(0+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<9))+(0+(layer_in_buffer[6]<<1)+(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<12))+(0-(layer_in_buffer[7]<<4)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<11)+(layer_in_buffer[7]<<12))-(0+(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<7)+(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<12))-(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<3)+(layer_in_buffer[9]<<6)+(layer_in_buffer[9]<<10))+(0+(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<3)-(layer_in_buffer[10]<<5)-(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<11))-(0-(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<6)-(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<11)+(layer_in_buffer[11]<<12))-(0-(layer_in_buffer[12]<<3)+(layer_in_buffer[12]<<8)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<11))-(0-(layer_in_buffer[13]<<3)-(layer_in_buffer[13]<<5)-(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<11)+(layer_in_buffer[13]<<12))-(0-(layer_in_buffer[14]<<1)+(layer_in_buffer[14]<<7)+(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<14))-(0+(layer_in_buffer[15]<<4)-(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<12))-(0+(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<4)+(layer_in_buffer[16]<<5)+(layer_in_buffer[16]<<11)+(layer_in_buffer[16]<<13))+(0+(layer_in_buffer[17]<<0)+(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<9))+(0+(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<6)+(layer_in_buffer[18]<<9))+(0-(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<4)-(layer_in_buffer[19]<<6)+(layer_in_buffer[19]<<10)+(layer_in_buffer[19]<<11))-(0+(layer_in_buffer[20]<<2)-(layer_in_buffer[20]<<5)-(layer_in_buffer[20]<<7)-(layer_in_buffer[20]<<9)+(layer_in_buffer[20]<<12)+(layer_in_buffer[20]<<13))+(0+(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<2)-(layer_in_buffer[21]<<5)+(layer_in_buffer[21]<<8)+(layer_in_buffer[21]<<10))+(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<1)-(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<9)+(layer_in_buffer[22]<<10))+(0+(layer_in_buffer[23]<<0)+(layer_in_buffer[23]<<3)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<8)+(layer_in_buffer[23]<<10)+(layer_in_buffer[23]<<13))+(0+(layer_in_buffer[24]<<1)+(layer_in_buffer[24]<<2)+(layer_in_buffer[24]<<5)+(layer_in_buffer[24]<<7))+(0+(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<1)-(layer_in_buffer[25]<<4)-(layer_in_buffer[25]<<6)-(layer_in_buffer[25]<<8)+(layer_in_buffer[25]<<10)+(layer_in_buffer[25]<<11))-(0+(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<2)+(layer_in_buffer[26]<<5)+(layer_in_buffer[26]<<6)-(layer_in_buffer[26]<<9)+(layer_in_buffer[26]<<12)+(layer_in_buffer[26]<<13))-(0-(layer_in_buffer[27]<<1)+(layer_in_buffer[27]<<5)+(layer_in_buffer[27]<<6)+(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<13))+(0+(layer_in_buffer[28]<<2)-(layer_in_buffer[28]<<5)+(layer_in_buffer[28]<<10))-(0+(layer_in_buffer[30]<<3)+(layer_in_buffer[30]<<4)+(layer_in_buffer[30]<<7)+(layer_in_buffer[30]<<9))-(0-(layer_in_buffer[31]<<0)+(layer_in_buffer[31]<<3)+(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<7)-(layer_in_buffer[31]<<9)+(layer_in_buffer[31]<<12))-(0-(layer_in_buffer[32]<<3)-(layer_in_buffer[32]<<6)+(layer_in_buffer[32]<<9)+(layer_in_buffer[32]<<13))-(0+(layer_in_buffer[33]<<1)+(layer_in_buffer[33]<<3)-(layer_in_buffer[33]<<5)-(layer_in_buffer[33]<<8)+(layer_in_buffer[33]<<12))-(0+(layer_in_buffer[34]<<0)+(layer_in_buffer[34]<<4)-(layer_in_buffer[34]<<6)+(layer_in_buffer[34]<<9)+(layer_in_buffer[34]<<14))+(0+(layer_in_buffer[35]<<3)+(layer_in_buffer[35]<<4)+(layer_in_buffer[35]<<7)+(layer_in_buffer[35]<<9))-(0+(layer_in_buffer[36]<<4)+(layer_in_buffer[36]<<5)+(layer_in_buffer[36]<<8)+(layer_in_buffer[36]<<10))+(0+(layer_in_buffer[37]<<1)+(layer_in_buffer[37]<<7)+(layer_in_buffer[37]<<8)+(layer_in_buffer[37]<<12))-(0+(layer_in_buffer[38]<<0)+(layer_in_buffer[38]<<2)+(layer_in_buffer[38]<<5)+(layer_in_buffer[38]<<7)+(layer_in_buffer[38]<<10)+(layer_in_buffer[38]<<11))+(0+(layer_in_buffer[39]<<1)-(layer_in_buffer[39]<<4)+(layer_in_buffer[39]<<9))+(0+(layer_in_buffer[40]<<2)+(layer_in_buffer[40]<<4)+(layer_in_buffer[40]<<8)+(layer_in_buffer[40]<<11))-(0+(layer_in_buffer[41]<<0)+(layer_in_buffer[41]<<1)-(layer_in_buffer[41]<<4)-(layer_in_buffer[41]<<6)-(layer_in_buffer[41]<<8)+(layer_in_buffer[41]<<10)+(layer_in_buffer[41]<<11))-(0+(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<2)+(layer_in_buffer[42]<<6)+(layer_in_buffer[42]<<9))-(0-(layer_in_buffer[43]<<1)+(layer_in_buffer[43]<<11)+(layer_in_buffer[43]<<12))+(0+(layer_in_buffer[44]<<0)-(layer_in_buffer[44]<<2)-(layer_in_buffer[44]<<5)+(layer_in_buffer[44]<<8)+(layer_in_buffer[44]<<10))+(0+(layer_in_buffer[45]<<0)+(layer_in_buffer[45]<<1)-(layer_in_buffer[45]<<4)-(layer_in_buffer[45]<<7)+(layer_in_buffer[45]<<13))+(0+(layer_in_buffer[46]<<0)+(layer_in_buffer[46]<<3)-(layer_in_buffer[46]<<5)-(layer_in_buffer[46]<<8)-(layer_in_buffer[46]<<10)+(layer_in_buffer[46]<<13))+(0+(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<5)+(layer_in_buffer[47]<<7)+(layer_in_buffer[47]<<11)+(layer_in_buffer[47]<<12))+(0-(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<4)-(layer_in_buffer[48]<<6)-(layer_in_buffer[48]<<8)+(layer_in_buffer[48]<<11))-(0-(layer_in_buffer[49]<<1)-(layer_in_buffer[49]<<3)-(layer_in_buffer[49]<<5)+(layer_in_buffer[49]<<9)+(layer_in_buffer[49]<<10))+(0-(layer_in_buffer[50]<<1)-(layer_in_buffer[50]<<3)+(layer_in_buffer[50]<<6)+(layer_in_buffer[50]<<12))-(0-(layer_in_buffer[51]<<6)+(layer_in_buffer[51]<<11)+(layer_in_buffer[51]<<13)+(layer_in_buffer[51]<<14))-(0+(layer_in_buffer[52]<<1)+(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<5)+(layer_in_buffer[52]<<7))-(0-(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<7)+(layer_in_buffer[53]<<9)+(layer_in_buffer[53]<<10))+(0+(layer_in_buffer[54]<<3)-(layer_in_buffer[54]<<6)+(layer_in_buffer[54]<<11))+(0+(layer_in_buffer[55]<<0)+(layer_in_buffer[55]<<2)+(layer_in_buffer[55]<<5)+(layer_in_buffer[55]<<7)+(layer_in_buffer[55]<<10)+(layer_in_buffer[55]<<11))+(0+(layer_in_buffer[56]<<6)+(layer_in_buffer[56]<<7)+(layer_in_buffer[56]<<10)+(layer_in_buffer[56]<<12))-(0+(layer_in_buffer[58]<<0)+(layer_in_buffer[58]<<6)+(layer_in_buffer[58]<<7)+(layer_in_buffer[58]<<11))-(0+(layer_in_buffer[59]<<0)+(layer_in_buffer[59]<<1)-(layer_in_buffer[59]<<6)+(layer_in_buffer[59]<<10)+(layer_in_buffer[59]<<14))+(0+(layer_in_buffer[60]<<0)-(layer_in_buffer[60]<<2)-(layer_in_buffer[60]<<5)+(layer_in_buffer[60]<<8)+(layer_in_buffer[60]<<10))+(0+(layer_in_buffer[61]<<1)+(layer_in_buffer[61]<<2)+(layer_in_buffer[61]<<5)+(layer_in_buffer[61]<<7))+(0-(layer_in_buffer[62]<<0)-(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<7)+(layer_in_buffer[62]<<9)+(layer_in_buffer[62]<<12))-(0+(layer_in_buffer[63]<<2)-(layer_in_buffer[63]<<5)+(layer_in_buffer[63]<<10));
wire [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0-(0+(layer_in_buffer[0]<<1)+(layer_in_buffer[0]<<2)-(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<11))+(0+(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<4)+(layer_in_buffer[1]<<7)+(layer_in_buffer[1]<<9)+(layer_in_buffer[1]<<12)+(layer_in_buffer[1]<<13))+(0+(layer_in_buffer[2]<<4)+(layer_in_buffer[2]<<5)-(layer_in_buffer[2]<<11)+(layer_in_buffer[2]<<13)+(layer_in_buffer[2]<<14))-(0-(layer_in_buffer[3]<<2)-(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<7)+(layer_in_buffer[3]<<13))+(0+(layer_in_buffer[4]<<1)+(layer_in_buffer[4]<<3)+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<10)+(layer_in_buffer[4]<<12))+(0+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<3)-(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<11)+(layer_in_buffer[5]<<12))+(0+(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<1)-(layer_in_buffer[6]<<5)+(layer_in_buffer[6]<<12))-(0+(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<2)-(layer_in_buffer[7]<<5)-(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<10)+(layer_in_buffer[7]<<11)+(layer_in_buffer[7]<<14))-(0+(layer_in_buffer[8]<<2)-(layer_in_buffer[8]<<4)-(layer_in_buffer[8]<<7)+(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<12))+(0+(layer_in_buffer[9]<<0)+(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<4)+(layer_in_buffer[9]<<6))-(0+(layer_in_buffer[10]<<3)+(layer_in_buffer[10]<<6)+(layer_in_buffer[10]<<8)+(layer_in_buffer[10]<<12)+(layer_in_buffer[10]<<13))+(0+(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<4)-(layer_in_buffer[11]<<6)+(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<13))+(0+(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<2)-(layer_in_buffer[12]<<4)-(layer_in_buffer[12]<<7)+(layer_in_buffer[12]<<11))-(0-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<12)+(layer_in_buffer[13]<<13))-(0-(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<3)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<13))-(0+(layer_in_buffer[15]<<1)+(layer_in_buffer[15]<<2)-(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<10)+(layer_in_buffer[15]<<11))-(0+(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<6)+(layer_in_buffer[16]<<7)-(layer_in_buffer[16]<<11)+(layer_in_buffer[16]<<14))-(0+(layer_in_buffer[17]<<3)+(layer_in_buffer[17]<<4)+(layer_in_buffer[17]<<7)+(layer_in_buffer[17]<<9))-(0+(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<4)+(layer_in_buffer[18]<<5)-(layer_in_buffer[18]<<10)+(layer_in_buffer[18]<<13))-(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<4)-(layer_in_buffer[19]<<6)+(layer_in_buffer[19]<<11)+(layer_in_buffer[19]<<12))-(0-(layer_in_buffer[20]<<2)-(layer_in_buffer[20]<<4)-(layer_in_buffer[20]<<6)+(layer_in_buffer[20]<<10)+(layer_in_buffer[20]<<11))-(0+(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<3)+(layer_in_buffer[21]<<10)+(layer_in_buffer[21]<<12)+(layer_in_buffer[21]<<14))-(0+(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<3)+(layer_in_buffer[22]<<8))-(0+(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<2)-(layer_in_buffer[23]<<5)-(layer_in_buffer[23]<<11)+(layer_in_buffer[23]<<13)+(layer_in_buffer[23]<<14))+(0+(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<4)+(layer_in_buffer[24]<<7)+(layer_in_buffer[24]<<9))+(0+(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<2)+(layer_in_buffer[26]<<5)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<8)+(layer_in_buffer[26]<<11)+(layer_in_buffer[26]<<12))-(0-(layer_in_buffer[27]<<1)-(layer_in_buffer[27]<<3)-(layer_in_buffer[27]<<5)+(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<10))-(0+(layer_in_buffer[28]<<4)+(layer_in_buffer[28]<<5)+(layer_in_buffer[28]<<8)+(layer_in_buffer[28]<<10))+(0-(layer_in_buffer[29]<<2)-(layer_in_buffer[29]<<5)+(layer_in_buffer[29]<<8)+(layer_in_buffer[29]<<12))-(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<4)+(layer_in_buffer[30]<<9)+(layer_in_buffer[30]<<10)+(layer_in_buffer[30]<<13))-(0-(layer_in_buffer[31]<<1)+(layer_in_buffer[31]<<5)+(layer_in_buffer[31]<<6)+(layer_in_buffer[31]<<9)+(layer_in_buffer[31]<<13))-(0+(layer_in_buffer[32]<<1)+(layer_in_buffer[32]<<3)+(layer_in_buffer[32]<<7)+(layer_in_buffer[32]<<10))+(0-(layer_in_buffer[33]<<2)-(layer_in_buffer[33]<<5)+(layer_in_buffer[33]<<8)+(layer_in_buffer[33]<<12))-(0+(layer_in_buffer[34]<<0)+(layer_in_buffer[34]<<2)+(layer_in_buffer[34]<<5)+(layer_in_buffer[34]<<7)+(layer_in_buffer[34]<<10)+(layer_in_buffer[34]<<11))+(0+(layer_in_buffer[35]<<0)-(layer_in_buffer[35]<<2)-(layer_in_buffer[35]<<5)+(layer_in_buffer[35]<<8)+(layer_in_buffer[35]<<10))-(0+(layer_in_buffer[36]<<0)-(layer_in_buffer[36]<<3)+(layer_in_buffer[36]<<7)+(layer_in_buffer[36]<<9)+(layer_in_buffer[36]<<11)+(layer_in_buffer[36]<<13))+(0+(layer_in_buffer[37]<<1)+(layer_in_buffer[37]<<3)+(layer_in_buffer[37]<<4)+(layer_in_buffer[37]<<10)+(layer_in_buffer[37]<<12))+(0-(layer_in_buffer[38]<<0)-(layer_in_buffer[38]<<2)-(layer_in_buffer[38]<<5)+(layer_in_buffer[38]<<8)-(layer_in_buffer[38]<<10)+(layer_in_buffer[38]<<13))-(0+(layer_in_buffer[39]<<4)-(layer_in_buffer[39]<<6)-(layer_in_buffer[39]<<9)+(layer_in_buffer[39]<<12)+(layer_in_buffer[39]<<14))+(0+(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<4)-(layer_in_buffer[40]<<9)+(layer_in_buffer[40]<<12))+(0-(layer_in_buffer[41]<<0)+(layer_in_buffer[41]<<4)-(layer_in_buffer[41]<<7)-(layer_in_buffer[41]<<10)+(layer_in_buffer[41]<<13))-(0+(layer_in_buffer[42]<<1)+(layer_in_buffer[42]<<2)+(layer_in_buffer[42]<<5)+(layer_in_buffer[42]<<7))-(0-(layer_in_buffer[43]<<2)-(layer_in_buffer[43]<<4)+(layer_in_buffer[43]<<9)+(layer_in_buffer[43]<<11)+(layer_in_buffer[43]<<14))-(0-(layer_in_buffer[44]<<0)-(layer_in_buffer[44]<<3)+(layer_in_buffer[44]<<6)+(layer_in_buffer[44]<<10))+(0-(layer_in_buffer[45]<<0)+(layer_in_buffer[45]<<5)-(layer_in_buffer[45]<<8)-(layer_in_buffer[45]<<10)+(layer_in_buffer[45]<<12)+(layer_in_buffer[45]<<13))-(0-(layer_in_buffer[46]<<0)+(layer_in_buffer[46]<<3)-(layer_in_buffer[46]<<5)+(layer_in_buffer[46]<<7)+(layer_in_buffer[46]<<8)+(layer_in_buffer[46]<<11))-(0+(layer_in_buffer[47]<<1)+(layer_in_buffer[47]<<4)+(layer_in_buffer[47]<<8)+(layer_in_buffer[47]<<13))-(0+(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<1)+(layer_in_buffer[48]<<4)+(layer_in_buffer[48]<<8)+(layer_in_buffer[48]<<10)+(layer_in_buffer[48]<<12))+(0+(layer_in_buffer[49]<<1)+(layer_in_buffer[49]<<3)+(layer_in_buffer[49]<<5)+(layer_in_buffer[49]<<8)+(layer_in_buffer[49]<<10)+(layer_in_buffer[49]<<11)+(layer_in_buffer[49]<<14))+(0+(layer_in_buffer[51]<<2)-(layer_in_buffer[51]<<4)-(layer_in_buffer[51]<<7)+(layer_in_buffer[51]<<10)+(layer_in_buffer[51]<<12))-(0+(layer_in_buffer[52]<<0)+(layer_in_buffer[52]<<2)+(layer_in_buffer[52]<<5)+(layer_in_buffer[52]<<7)+(layer_in_buffer[52]<<10)+(layer_in_buffer[52]<<11))-(0+(layer_in_buffer[53]<<0)-(layer_in_buffer[53]<<7)-(layer_in_buffer[53]<<9)+(layer_in_buffer[53]<<13))-(0-(layer_in_buffer[54]<<0)+(layer_in_buffer[54]<<3)-(layer_in_buffer[54]<<5)+(layer_in_buffer[54]<<7)+(layer_in_buffer[54]<<8)+(layer_in_buffer[54]<<11))+(0+(layer_in_buffer[55]<<3)+(layer_in_buffer[55]<<4)+(layer_in_buffer[55]<<7)+(layer_in_buffer[55]<<9))-(0+(layer_in_buffer[56]<<1)+(layer_in_buffer[56]<<2)-(layer_in_buffer[56]<<6)+(layer_in_buffer[56]<<13))+(0+(layer_in_buffer[57]<<0)-(layer_in_buffer[57]<<2)-(layer_in_buffer[57]<<5)+(layer_in_buffer[57]<<8)+(layer_in_buffer[57]<<10))+(0+(layer_in_buffer[58]<<0)+(layer_in_buffer[58]<<3)+(layer_in_buffer[58]<<9)-(layer_in_buffer[58]<<11)+(layer_in_buffer[58]<<14))-(0+(layer_in_buffer[59]<<0)-(layer_in_buffer[59]<<2)-(layer_in_buffer[59]<<4)-(layer_in_buffer[59]<<9)+(layer_in_buffer[59]<<14))-(0+(layer_in_buffer[60]<<1)+(layer_in_buffer[60]<<3)+(layer_in_buffer[60]<<4)+(layer_in_buffer[60]<<10)+(layer_in_buffer[60]<<12))-(0+(layer_in_buffer[61]<<3)+(layer_in_buffer[61]<<4)+(layer_in_buffer[61]<<7)+(layer_in_buffer[61]<<9))-(0+(layer_in_buffer[62]<<3)+(layer_in_buffer[62]<<5)+(layer_in_buffer[62]<<9)+(layer_in_buffer[62]<<12))-(0+(layer_in_buffer[63]<<2)-(layer_in_buffer[63]<<5)+(layer_in_buffer[63]<<10));
wire [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0-(0+(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<6)-(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<11)+(layer_in_buffer[0]<<14))-(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<11))-(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)-(layer_in_buffer[2]<<4)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<9))+(0+(layer_in_buffer[3]<<4)-(layer_in_buffer[3]<<7)+(layer_in_buffer[3]<<12))-(0+(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<4)+(layer_in_buffer[4]<<6)+(layer_in_buffer[4]<<11)+(layer_in_buffer[4]<<12))-(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<1)-(layer_in_buffer[5]<<5)+(layer_in_buffer[5]<<12))+(0+(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<7)+(layer_in_buffer[6]<<9)+(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<13))+(0+(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<3)+(layer_in_buffer[7]<<6)+(layer_in_buffer[7]<<8))+(0-(layer_in_buffer[8]<<1)+(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<9))+(0+(layer_in_buffer[9]<<0)+(layer_in_buffer[9]<<4)-(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<10))+(0-(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<3)+(layer_in_buffer[10]<<4)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<9)+(layer_in_buffer[10]<<11)+(layer_in_buffer[10]<<12))+(0+(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<2)-(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<10))+(0+(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<2)+(layer_in_buffer[12]<<6)+(layer_in_buffer[12]<<9))-(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<2)-(layer_in_buffer[13]<<4)-(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<11))-(0+(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<6)+(layer_in_buffer[14]<<7)-(layer_in_buffer[14]<<11)+(layer_in_buffer[14]<<14))+(0+(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<5)+(layer_in_buffer[15]<<9)+(layer_in_buffer[15]<<10))-(0+(layer_in_buffer[16]<<0)+(layer_in_buffer[16]<<5)+(layer_in_buffer[16]<<8)+(layer_in_buffer[16]<<9)+(layer_in_buffer[16]<<12))-(0-(layer_in_buffer[17]<<0)+(layer_in_buffer[17]<<5)+(layer_in_buffer[17]<<7)+(layer_in_buffer[17]<<8))+(0-(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<5)+(layer_in_buffer[18]<<7)+(layer_in_buffer[18]<<8))+(0-(layer_in_buffer[19]<<0)+(layer_in_buffer[19]<<4)-(layer_in_buffer[19]<<6)-(layer_in_buffer[19]<<8)+(layer_in_buffer[19]<<11))+(0-(layer_in_buffer[20]<<1)+(layer_in_buffer[20]<<5)-(layer_in_buffer[20]<<7)-(layer_in_buffer[20]<<9)+(layer_in_buffer[20]<<12))+(0-(layer_in_buffer[21]<<1)-(layer_in_buffer[21]<<3)-(layer_in_buffer[21]<<5)+(layer_in_buffer[21]<<9)+(layer_in_buffer[21]<<10))+(0-(layer_in_buffer[22]<<1)-(layer_in_buffer[22]<<4)+(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<11))-(0-(layer_in_buffer[23]<<2)+(layer_in_buffer[23]<<5)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<9)-(layer_in_buffer[23]<<11)+(layer_in_buffer[23]<<14))-(0+(layer_in_buffer[24]<<1)+(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<7)+(layer_in_buffer[24]<<10))+(0+(layer_in_buffer[25]<<2)-(layer_in_buffer[25]<<5)+(layer_in_buffer[25]<<10))-(0-(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<3)+(layer_in_buffer[26]<<8)+(layer_in_buffer[26]<<11)+(layer_in_buffer[26]<<12))+(0+(layer_in_buffer[27]<<0)+(layer_in_buffer[27]<<4)+(layer_in_buffer[27]<<6)+(layer_in_buffer[27]<<11)+(layer_in_buffer[27]<<12))+(0+(layer_in_buffer[28]<<1)+(layer_in_buffer[28]<<3)+(layer_in_buffer[28]<<4)+(layer_in_buffer[28]<<10)+(layer_in_buffer[28]<<12))-(0+(layer_in_buffer[29]<<1)-(layer_in_buffer[29]<<4)+(layer_in_buffer[29]<<9))-(0+(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<1)-(layer_in_buffer[30]<<5)+(layer_in_buffer[30]<<12))+(0-(layer_in_buffer[31]<<0)+(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<3)+(layer_in_buffer[31]<<6)+(layer_in_buffer[31]<<8)+(layer_in_buffer[31]<<10)+(layer_in_buffer[31]<<11))-(0+(layer_in_buffer[32]<<2)+(layer_in_buffer[32]<<6)-(layer_in_buffer[32]<<9)+(layer_in_buffer[32]<<12))-(0+(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<2)-(layer_in_buffer[33]<<5)+(layer_in_buffer[33]<<8)+(layer_in_buffer[33]<<10))-(0+(layer_in_buffer[34]<<2)+(layer_in_buffer[34]<<8)+(layer_in_buffer[34]<<9)+(layer_in_buffer[34]<<13))-(0+(layer_in_buffer[35]<<0)+(layer_in_buffer[35]<<2)+(layer_in_buffer[35]<<6)+(layer_in_buffer[35]<<9))-(0+(layer_in_buffer[36]<<0)+(layer_in_buffer[36]<<2)+(layer_in_buffer[36]<<5)+(layer_in_buffer[36]<<7)+(layer_in_buffer[36]<<10)+(layer_in_buffer[36]<<11))-(0+(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<2)+(layer_in_buffer[37]<<5)+(layer_in_buffer[37]<<6)-(layer_in_buffer[37]<<9)+(layer_in_buffer[37]<<12)+(layer_in_buffer[37]<<13))+(0+(layer_in_buffer[38]<<0)+(layer_in_buffer[38]<<2)-(layer_in_buffer[38]<<4)-(layer_in_buffer[38]<<7)+(layer_in_buffer[38]<<11))+(0+(layer_in_buffer[39]<<2)-(layer_in_buffer[39]<<5)+(layer_in_buffer[39]<<10))-(0-(layer_in_buffer[40]<<1)+(layer_in_buffer[40]<<6)+(layer_in_buffer[40]<<8)+(layer_in_buffer[40]<<9))+(0+(layer_in_buffer[41]<<0)+(layer_in_buffer[41]<<4)-(layer_in_buffer[41]<<7)+(layer_in_buffer[41]<<10))+(0+(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<3)+(layer_in_buffer[42]<<5)+(layer_in_buffer[42]<<9)+(layer_in_buffer[42]<<10))+(0-(layer_in_buffer[43]<<0)+(layer_in_buffer[43]<<2)+(layer_in_buffer[43]<<3)+(layer_in_buffer[43]<<6)+(layer_in_buffer[43]<<8)+(layer_in_buffer[43]<<10)+(layer_in_buffer[43]<<11))-(0+(layer_in_buffer[44]<<0)-(layer_in_buffer[44]<<3)+(layer_in_buffer[44]<<8))+(0+(layer_in_buffer[45]<<5)+(layer_in_buffer[45]<<6)+(layer_in_buffer[45]<<9)+(layer_in_buffer[45]<<11))-(0-(layer_in_buffer[46]<<0)+(layer_in_buffer[46]<<4)+(layer_in_buffer[46]<<6)+(layer_in_buffer[46]<<12)+(layer_in_buffer[46]<<13))-(0+(layer_in_buffer[47]<<0)+(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<5)-(layer_in_buffer[47]<<9)-(layer_in_buffer[47]<<11)+(layer_in_buffer[47]<<14))+(0-(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<3)-(layer_in_buffer[48]<<5)+(layer_in_buffer[48]<<7)+(layer_in_buffer[48]<<8)+(layer_in_buffer[48]<<11))-(0-(layer_in_buffer[49]<<1)-(layer_in_buffer[49]<<4)+(layer_in_buffer[49]<<7)+(layer_in_buffer[49]<<11))+(0+(layer_in_buffer[50]<<0)-(layer_in_buffer[50]<<2)+(layer_in_buffer[50]<<6)-(layer_in_buffer[50]<<8)+(layer_in_buffer[50]<<12))-(0-(layer_in_buffer[51]<<0)+(layer_in_buffer[51]<<3)+(layer_in_buffer[51]<<5)+(layer_in_buffer[51]<<8)-(layer_in_buffer[51]<<12)+(layer_in_buffer[51]<<15))+(0+(layer_in_buffer[52]<<1)+(layer_in_buffer[52]<<3)+(layer_in_buffer[52]<<7)+(layer_in_buffer[52]<<10))-(0+(layer_in_buffer[53]<<0)+(layer_in_buffer[53]<<2)+(layer_in_buffer[53]<<6)+(layer_in_buffer[53]<<9))+(0-(layer_in_buffer[54]<<1)+(layer_in_buffer[54]<<6)+(layer_in_buffer[54]<<8)+(layer_in_buffer[54]<<9))-(0+(layer_in_buffer[55]<<4)-(layer_in_buffer[55]<<7)+(layer_in_buffer[55]<<12))+(0-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<7)+(layer_in_buffer[56]<<9)+(layer_in_buffer[56]<<10))-(0-(layer_in_buffer[57]<<3)+(layer_in_buffer[57]<<8)+(layer_in_buffer[57]<<10)+(layer_in_buffer[57]<<11))+(0+(layer_in_buffer[58]<<1)+(layer_in_buffer[58]<<3)+(layer_in_buffer[58]<<6)+(layer_in_buffer[58]<<8)+(layer_in_buffer[58]<<11)+(layer_in_buffer[58]<<12))+(0+(layer_in_buffer[59]<<7)+(layer_in_buffer[59]<<8)+(layer_in_buffer[59]<<11)+(layer_in_buffer[59]<<13))+(0+(layer_in_buffer[60]<<0)+(layer_in_buffer[60]<<3)+(layer_in_buffer[60]<<5)+(layer_in_buffer[60]<<9)+(layer_in_buffer[60]<<10))+(0+(layer_in_buffer[61]<<0)+(layer_in_buffer[61]<<2)+(layer_in_buffer[61]<<3)+(layer_in_buffer[61]<<9)+(layer_in_buffer[61]<<11))+(0+(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<3)+(layer_in_buffer[62]<<6)+(layer_in_buffer[62]<<8))-(0+(layer_in_buffer[63]<<0)+(layer_in_buffer[63]<<4)-(layer_in_buffer[63]<<7)+(layer_in_buffer[63]<<10));
wire [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0-(0+(layer_in_buffer[0]<<1)-(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<6)+(layer_in_buffer[0]<<7)-(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<13)+(layer_in_buffer[0]<<14))+(0-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<6)-(layer_in_buffer[1]<<8)-(layer_in_buffer[1]<<10)+(layer_in_buffer[1]<<13))-(0+(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<1)-(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<12))+(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<1)+(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<12))-(0-(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<2)+(layer_in_buffer[4]<<6)-(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<11)+(layer_in_buffer[4]<<13))+(0-(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<3)+(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<7)-(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<12))-(0+(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<2)+(layer_in_buffer[6]<<3)-(layer_in_buffer[6]<<6)-(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<13))-(0+(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<13))-(0+(layer_in_buffer[8]<<4)+(layer_in_buffer[8]<<5)+(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<10))+(0-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<7)+(layer_in_buffer[9]<<9)+(layer_in_buffer[9]<<10))-(0-(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)-(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<8)-(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<13))+(0+(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<5)+(layer_in_buffer[11]<<8)+(layer_in_buffer[11]<<10))-(0-(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<11))+(0+(layer_in_buffer[13]<<1)+(layer_in_buffer[13]<<2)-(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<11))+(0+(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<4)-(layer_in_buffer[14]<<7)-(layer_in_buffer[14]<<11)+(layer_in_buffer[14]<<14))-(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<10))+(0-(layer_in_buffer[16]<<4)-(layer_in_buffer[16]<<6)-(layer_in_buffer[16]<<8)+(layer_in_buffer[16]<<12)+(layer_in_buffer[16]<<13))+(0+(layer_in_buffer[17]<<1)-(layer_in_buffer[17]<<3)-(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<9)+(layer_in_buffer[17]<<11))+(0+(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<4)+(layer_in_buffer[18]<<6)+(layer_in_buffer[18]<<11)+(layer_in_buffer[18]<<12))-(0-(layer_in_buffer[19]<<0)+(layer_in_buffer[19]<<4)-(layer_in_buffer[19]<<7)-(layer_in_buffer[19]<<10)+(layer_in_buffer[19]<<13))+(0+(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<1)+(layer_in_buffer[20]<<4)+(layer_in_buffer[20]<<8)+(layer_in_buffer[20]<<10)+(layer_in_buffer[20]<<12))-(0+(layer_in_buffer[21]<<3)-(layer_in_buffer[21]<<6)+(layer_in_buffer[21]<<11))+(0-(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<11))-(0+(layer_in_buffer[23]<<0)+(layer_in_buffer[23]<<2)-(layer_in_buffer[23]<<5)+(layer_in_buffer[23]<<7)+(layer_in_buffer[23]<<8)+(layer_in_buffer[23]<<13))+(0+(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<3)+(layer_in_buffer[25]<<5)+(layer_in_buffer[25]<<9)+(layer_in_buffer[25]<<10))-(0+(layer_in_buffer[26]<<0)+(layer_in_buffer[26]<<2)-(layer_in_buffer[26]<<4)-(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<11))-(0+(layer_in_buffer[27]<<1)-(layer_in_buffer[27]<<4)-(layer_in_buffer[27]<<6)-(layer_in_buffer[27]<<8)+(layer_in_buffer[27]<<11)+(layer_in_buffer[27]<<12))+(0-(layer_in_buffer[28]<<0)+(layer_in_buffer[28]<<10)+(layer_in_buffer[28]<<11))-(0+(layer_in_buffer[29]<<3)+(layer_in_buffer[29]<<4)+(layer_in_buffer[29]<<7)+(layer_in_buffer[29]<<9))+(0+(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<1)-(layer_in_buffer[30]<<7)+(layer_in_buffer[30]<<9)+(layer_in_buffer[30]<<10))-(0-(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<9)+(layer_in_buffer[31]<<11)+(layer_in_buffer[31]<<12))+(0+(layer_in_buffer[32]<<2)-(layer_in_buffer[32]<<5)+(layer_in_buffer[32]<<10))-(0-(layer_in_buffer[33]<<0)+(layer_in_buffer[33]<<4)+(layer_in_buffer[33]<<5)+(layer_in_buffer[33]<<8)+(layer_in_buffer[33]<<12))+(0+(layer_in_buffer[34]<<0)+(layer_in_buffer[34]<<3)-(layer_in_buffer[34]<<5)-(layer_in_buffer[34]<<8)-(layer_in_buffer[34]<<10)+(layer_in_buffer[34]<<13))+(0-(layer_in_buffer[36]<<0)+(layer_in_buffer[36]<<5)+(layer_in_buffer[36]<<7)+(layer_in_buffer[36]<<8))+(0+(layer_in_buffer[37]<<4)+(layer_in_buffer[37]<<5)+(layer_in_buffer[37]<<8)+(layer_in_buffer[37]<<10))+(0+(layer_in_buffer[38]<<3)+(layer_in_buffer[38]<<4)+(layer_in_buffer[38]<<7)+(layer_in_buffer[38]<<9))-(0+(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<4)+(layer_in_buffer[39]<<8)+(layer_in_buffer[39]<<11))+(0+(layer_in_buffer[40]<<1)-(layer_in_buffer[40]<<4)+(layer_in_buffer[40]<<9))-(0+(layer_in_buffer[41]<<6)+(layer_in_buffer[41]<<7)+(layer_in_buffer[41]<<10)+(layer_in_buffer[41]<<12))+(0+(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<1)-(layer_in_buffer[42]<<7)+(layer_in_buffer[42]<<9)+(layer_in_buffer[42]<<10))-(0-(layer_in_buffer[43]<<0)-(layer_in_buffer[43]<<3)+(layer_in_buffer[43]<<6)+(layer_in_buffer[43]<<10))+(0-(layer_in_buffer[44]<<2)-(layer_in_buffer[44]<<4)-(layer_in_buffer[44]<<6)+(layer_in_buffer[44]<<10)+(layer_in_buffer[44]<<11))-(0+(layer_in_buffer[45]<<1)-(layer_in_buffer[45]<<3)+(layer_in_buffer[45]<<6)+(layer_in_buffer[45]<<8)+(layer_in_buffer[45]<<9)+(layer_in_buffer[45]<<12)+(layer_in_buffer[45]<<13))-(0-(layer_in_buffer[46]<<2)+(layer_in_buffer[46]<<6)-(layer_in_buffer[46]<<8)-(layer_in_buffer[46]<<10)+(layer_in_buffer[46]<<13))-(0-(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<2)-(layer_in_buffer[47]<<4)-(layer_in_buffer[47]<<6)+(layer_in_buffer[47]<<11)+(layer_in_buffer[47]<<12))-(0-(layer_in_buffer[48]<<1)+(layer_in_buffer[48]<<7)+(layer_in_buffer[48]<<8)+(layer_in_buffer[48]<<14))-(0-(layer_in_buffer[49]<<0)+(layer_in_buffer[49]<<10)+(layer_in_buffer[49]<<11))-(0-(layer_in_buffer[50]<<0)-(layer_in_buffer[50]<<2)-(layer_in_buffer[50]<<4)+(layer_in_buffer[50]<<8)+(layer_in_buffer[50]<<9))+(0-(layer_in_buffer[51]<<0)+(layer_in_buffer[51]<<3)-(layer_in_buffer[51]<<5)+(layer_in_buffer[51]<<7)+(layer_in_buffer[51]<<8)+(layer_in_buffer[51]<<11))+(0+(layer_in_buffer[52]<<1)+(layer_in_buffer[52]<<4)+(layer_in_buffer[52]<<6)+(layer_in_buffer[52]<<10)+(layer_in_buffer[52]<<11))+(0+(layer_in_buffer[54]<<2)-(layer_in_buffer[54]<<5)+(layer_in_buffer[54]<<10))-(0-(layer_in_buffer[55]<<0)+(layer_in_buffer[55]<<4)-(layer_in_buffer[55]<<7)-(layer_in_buffer[55]<<10)+(layer_in_buffer[55]<<13))-(0-(layer_in_buffer[56]<<0)+(layer_in_buffer[56]<<10)+(layer_in_buffer[56]<<11))+(0+(layer_in_buffer[57]<<0)+(layer_in_buffer[57]<<1)-(layer_in_buffer[57]<<8)+(layer_in_buffer[57]<<12)+(layer_in_buffer[57]<<13))-(0+(layer_in_buffer[58]<<0)+(layer_in_buffer[58]<<6)+(layer_in_buffer[58]<<7)+(layer_in_buffer[58]<<11))-(0+(layer_in_buffer[59]<<1)+(layer_in_buffer[59]<<6)+(layer_in_buffer[59]<<8)-(layer_in_buffer[59]<<11)+(layer_in_buffer[59]<<15))+(0+(layer_in_buffer[60]<<0)+(layer_in_buffer[60]<<1)+(layer_in_buffer[60]<<4)+(layer_in_buffer[60]<<6))+(0-(layer_in_buffer[61]<<0)+(layer_in_buffer[61]<<10)+(layer_in_buffer[61]<<11))+(0-(layer_in_buffer[62]<<1)-(layer_in_buffer[62]<<3)+(layer_in_buffer[62]<<6)+(layer_in_buffer[62]<<12))+(0+(layer_in_buffer[63]<<2)+(layer_in_buffer[63]<<3)+(layer_in_buffer[63]<<6)+(layer_in_buffer[63]<<8));
wire [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0-(0-(layer_in_buffer[0]<<1)+(layer_in_buffer[0]<<3)+(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<7)+(layer_in_buffer[0]<<9)+(layer_in_buffer[0]<<11)+(layer_in_buffer[0]<<12))+(0+(layer_in_buffer[1]<<1)+(layer_in_buffer[1]<<3)+(layer_in_buffer[1]<<6)+(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<12))-(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)-(layer_in_buffer[2]<<4)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<9))-(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6)+(layer_in_buffer[3]<<9))-(0+(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<4)-(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<11))-(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<4)-(layer_in_buffer[5]<<6)+(layer_in_buffer[5]<<9)+(layer_in_buffer[5]<<12))-(0-(layer_in_buffer[6]<<1)+(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<8)+(layer_in_buffer[6]<<12)+(layer_in_buffer[6]<<14))+(0-(layer_in_buffer[7]<<1)+(layer_in_buffer[7]<<4)+(layer_in_buffer[7]<<5)+(layer_in_buffer[7]<<8)-(layer_in_buffer[7]<<10)+(layer_in_buffer[7]<<13))+(0+(layer_in_buffer[8]<<1)+(layer_in_buffer[8]<<5)-(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<11))+(0-(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<2)+(layer_in_buffer[9]<<5)+(layer_in_buffer[9]<<11))-(0+(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<8)+(layer_in_buffer[10]<<11)+(layer_in_buffer[10]<<12))+(0-(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<3)-(layer_in_buffer[11]<<6)+(layer_in_buffer[11]<<10)+(layer_in_buffer[11]<<12))+(0+(layer_in_buffer[12]<<1)+(layer_in_buffer[12]<<2)-(layer_in_buffer[12]<<8)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<11))-(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<4)+(layer_in_buffer[13]<<5)-(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<13))-(0+(layer_in_buffer[14]<<2)+(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<5)+(layer_in_buffer[14]<<11)+(layer_in_buffer[14]<<13))+(0-(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<4)-(layer_in_buffer[15]<<6)-(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<11))+(0+(layer_in_buffer[16]<<0)+(layer_in_buffer[16]<<2)+(layer_in_buffer[16]<<5)+(layer_in_buffer[16]<<7)+(layer_in_buffer[16]<<10)+(layer_in_buffer[16]<<11))-(0+(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<3)+(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<8))-(0-(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<10)+(layer_in_buffer[18]<<11))+(0+(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<8)+(layer_in_buffer[19]<<10))-(0+(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<2)-(layer_in_buffer[20]<<4)-(layer_in_buffer[20]<<7)+(layer_in_buffer[20]<<11))-(0-(layer_in_buffer[21]<<0)+(layer_in_buffer[21]<<5)+(layer_in_buffer[21]<<6)-(layer_in_buffer[21]<<9)+(layer_in_buffer[21]<<11)+(layer_in_buffer[21]<<12))+(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<2)-(layer_in_buffer[22]<<4)-(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<11))-(0+(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<7)-(layer_in_buffer[23]<<9)+(layer_in_buffer[23]<<13))-(0+(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<4)+(layer_in_buffer[24]<<7)+(layer_in_buffer[24]<<9))-(0+(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<4)-(layer_in_buffer[25]<<7)+(layer_in_buffer[25]<<10))-(0-(layer_in_buffer[26]<<1)-(layer_in_buffer[26]<<4)+(layer_in_buffer[26]<<7)+(layer_in_buffer[26]<<11))+(0+(layer_in_buffer[27]<<1)-(layer_in_buffer[27]<<3)-(layer_in_buffer[27]<<6)+(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<11))-(0-(layer_in_buffer[28]<<0)+(layer_in_buffer[28]<<4)-(layer_in_buffer[28]<<6)-(layer_in_buffer[28]<<8)+(layer_in_buffer[28]<<11))+(0+(layer_in_buffer[29]<<3)-(layer_in_buffer[29]<<6)+(layer_in_buffer[29]<<11))-(0+(layer_in_buffer[30]<<5)-(layer_in_buffer[30]<<8)+(layer_in_buffer[30]<<13))+(0+(layer_in_buffer[31]<<2)+(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<8)+(layer_in_buffer[31]<<11))+(0+(layer_in_buffer[32]<<3)+(layer_in_buffer[32]<<4)+(layer_in_buffer[32]<<7)+(layer_in_buffer[32]<<9))-(0+(layer_in_buffer[33]<<0)+(layer_in_buffer[33]<<1)+(layer_in_buffer[33]<<4)+(layer_in_buffer[33]<<6))+(0-(layer_in_buffer[34]<<0)+(layer_in_buffer[34]<<3)+(layer_in_buffer[34]<<7)+(layer_in_buffer[34]<<11)+(layer_in_buffer[34]<<13))+(0+(layer_in_buffer[35]<<0)+(layer_in_buffer[35]<<4)-(layer_in_buffer[35]<<7)+(layer_in_buffer[35]<<10))+(0+(layer_in_buffer[36]<<0)+(layer_in_buffer[36]<<2)+(layer_in_buffer[36]<<3)+(layer_in_buffer[36]<<9)+(layer_in_buffer[36]<<11))-(0+(layer_in_buffer[37]<<1)+(layer_in_buffer[37]<<3)+(layer_in_buffer[37]<<7)+(layer_in_buffer[37]<<10))-(0-(layer_in_buffer[38]<<3)+(layer_in_buffer[38]<<8)+(layer_in_buffer[38]<<10)+(layer_in_buffer[38]<<11))+(0+(layer_in_buffer[39]<<0)+(layer_in_buffer[39]<<2)-(layer_in_buffer[39]<<4)-(layer_in_buffer[39]<<7)+(layer_in_buffer[39]<<11))-(0+(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<3)+(layer_in_buffer[40]<<8))-(0-(layer_in_buffer[41]<<0)+(layer_in_buffer[41]<<5)+(layer_in_buffer[41]<<6)-(layer_in_buffer[41]<<9)+(layer_in_buffer[41]<<11)+(layer_in_buffer[41]<<12))+(0+(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<1)-(layer_in_buffer[42]<<7)+(layer_in_buffer[42]<<9)+(layer_in_buffer[42]<<10))+(0+(layer_in_buffer[43]<<0)+(layer_in_buffer[43]<<1)+(layer_in_buffer[43]<<6)+(layer_in_buffer[43]<<9)+(layer_in_buffer[43]<<11)+(layer_in_buffer[43]<<12))+(0+(layer_in_buffer[44]<<1)+(layer_in_buffer[44]<<2)+(layer_in_buffer[44]<<5)+(layer_in_buffer[44]<<7))+(0+(layer_in_buffer[45]<<1)-(layer_in_buffer[45]<<3)-(layer_in_buffer[45]<<6)+(layer_in_buffer[45]<<9)+(layer_in_buffer[45]<<11))-(0-(layer_in_buffer[46]<<0)+(layer_in_buffer[46]<<10)+(layer_in_buffer[46]<<11))-(0+(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<4)+(layer_in_buffer[47]<<6)-(layer_in_buffer[47]<<8)+(layer_in_buffer[47]<<11)+(layer_in_buffer[47]<<14))-(0+(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<6)+(layer_in_buffer[48]<<7)+(layer_in_buffer[48]<<11))+(0+(layer_in_buffer[49]<<0)+(layer_in_buffer[49]<<2)+(layer_in_buffer[49]<<6)+(layer_in_buffer[49]<<9))-(0-(layer_in_buffer[50]<<1)+(layer_in_buffer[50]<<6)+(layer_in_buffer[50]<<8)+(layer_in_buffer[50]<<9))+(0+(layer_in_buffer[51]<<1)+(layer_in_buffer[51]<<7)+(layer_in_buffer[51]<<8)+(layer_in_buffer[51]<<12))+(0-(layer_in_buffer[52]<<1)-(layer_in_buffer[52]<<3)-(layer_in_buffer[52]<<5)+(layer_in_buffer[52]<<9)+(layer_in_buffer[52]<<10))-(0-(layer_in_buffer[53]<<0)+(layer_in_buffer[53]<<10)+(layer_in_buffer[53]<<11))+(0+(layer_in_buffer[54]<<3)-(layer_in_buffer[54]<<6)+(layer_in_buffer[54]<<11))-(0+(layer_in_buffer[55]<<0)-(layer_in_buffer[55]<<7)-(layer_in_buffer[55]<<9)+(layer_in_buffer[55]<<13))+(0+(layer_in_buffer[56]<<1)+(layer_in_buffer[56]<<3)+(layer_in_buffer[56]<<7)+(layer_in_buffer[56]<<10))-(0-(layer_in_buffer[57]<<0)+(layer_in_buffer[57]<<3)+(layer_in_buffer[57]<<9)+(layer_in_buffer[57]<<12)+(layer_in_buffer[57]<<14))-(0+(layer_in_buffer[58]<<0)-(layer_in_buffer[58]<<2)+(layer_in_buffer[58]<<6)-(layer_in_buffer[58]<<8)+(layer_in_buffer[58]<<12))+(0+(layer_in_buffer[59]<<2)+(layer_in_buffer[59]<<4)+(layer_in_buffer[59]<<5)+(layer_in_buffer[59]<<11)+(layer_in_buffer[59]<<13))+(0+(layer_in_buffer[60]<<2)-(layer_in_buffer[60]<<5)+(layer_in_buffer[60]<<10))+(0-(layer_in_buffer[61]<<1)-(layer_in_buffer[61]<<3)-(layer_in_buffer[61]<<5)+(layer_in_buffer[61]<<9)+(layer_in_buffer[61]<<10))-(0+(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<6)-(layer_in_buffer[62]<<9)+(layer_in_buffer[62]<<12))+(0+(layer_in_buffer[63]<<0)+(layer_in_buffer[63]<<1)+(layer_in_buffer[63]<<4)+(layer_in_buffer[63]<<6));
wire [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0+(0+(layer_in_buffer[0]<<0)+(layer_in_buffer[0]<<2)-(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<11)+(layer_in_buffer[0]<<12))+(0-(layer_in_buffer[1]<<2)+(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<6)+(layer_in_buffer[1]<<9)-(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<14))+(0-(layer_in_buffer[2]<<2)-(layer_in_buffer[2]<<4)+(layer_in_buffer[2]<<7)+(layer_in_buffer[2]<<13))-(0-(layer_in_buffer[3]<<4)+(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<11)+(layer_in_buffer[3]<<12))-(0+(layer_in_buffer[4]<<0)-(layer_in_buffer[4]<<3)+(layer_in_buffer[4]<<8))+(0+(layer_in_buffer[5]<<1)+(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<8)+(layer_in_buffer[5]<<12))-(0-(layer_in_buffer[6]<<1)+(layer_in_buffer[6]<<4)-(layer_in_buffer[6]<<7)+(layer_in_buffer[6]<<11)+(layer_in_buffer[6]<<13))+(0+(layer_in_buffer[7]<<2)+(layer_in_buffer[7]<<4)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<11))+(0+(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<3)-(layer_in_buffer[8]<<7)+(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<12)+(layer_in_buffer[8]<<13))-(0+(layer_in_buffer[9]<<0)-(layer_in_buffer[9]<<3)+(layer_in_buffer[9]<<8))+(0+(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<3)+(layer_in_buffer[10]<<6)+(layer_in_buffer[10]<<8))+(0+(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<2)+(layer_in_buffer[11]<<7)+(layer_in_buffer[11]<<10)+(layer_in_buffer[11]<<12)+(layer_in_buffer[11]<<13))-(0-(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)-(layer_in_buffer[12]<<5)+(layer_in_buffer[12]<<8)-(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<13))+(0-(layer_in_buffer[13]<<0)-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<7)+(layer_in_buffer[13]<<9)+(layer_in_buffer[13]<<12))-(0-(layer_in_buffer[14]<<3)+(layer_in_buffer[14]<<6)-(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<10)+(layer_in_buffer[14]<<11)+(layer_in_buffer[14]<<14))-(0+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<4)+(layer_in_buffer[15]<<7)+(layer_in_buffer[15]<<9))+(0-(layer_in_buffer[16]<<0)-(layer_in_buffer[16]<<4)+(layer_in_buffer[16]<<9)+(layer_in_buffer[16]<<10)+(layer_in_buffer[16]<<13))+(0-(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<2)-(layer_in_buffer[17]<<4)-(layer_in_buffer[17]<<6)+(layer_in_buffer[17]<<11)+(layer_in_buffer[17]<<12))-(0-(layer_in_buffer[18]<<0)+(layer_in_buffer[18]<<3)+(layer_in_buffer[18]<<5)-(layer_in_buffer[18]<<9)+(layer_in_buffer[18]<<13))+(0-(layer_in_buffer[19]<<1)-(layer_in_buffer[19]<<3)-(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<9)+(layer_in_buffer[19]<<10))+(0-(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<3)-(layer_in_buffer[20]<<5)+(layer_in_buffer[20]<<7)+(layer_in_buffer[20]<<8)+(layer_in_buffer[20]<<11))-(0+(layer_in_buffer[21]<<0)+(layer_in_buffer[21]<<2)+(layer_in_buffer[21]<<3)+(layer_in_buffer[21]<<9)+(layer_in_buffer[21]<<11))-(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<6)+(layer_in_buffer[22]<<9)+(layer_in_buffer[22]<<12)+(layer_in_buffer[22]<<13))+(0+(layer_in_buffer[23]<<1)-(layer_in_buffer[23]<<4)-(layer_in_buffer[23]<<6)-(layer_in_buffer[23]<<8)+(layer_in_buffer[23]<<11)+(layer_in_buffer[23]<<12))-(0+(layer_in_buffer[24]<<1)+(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<7)+(layer_in_buffer[24]<<10))-(0+(layer_in_buffer[25]<<0)-(layer_in_buffer[25]<<2)+(layer_in_buffer[25]<<6)-(layer_in_buffer[25]<<8)+(layer_in_buffer[25]<<12))+(0+(layer_in_buffer[26]<<5)+(layer_in_buffer[26]<<6)+(layer_in_buffer[26]<<9)+(layer_in_buffer[26]<<11))+(0+(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6)-(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<12))-(0+(layer_in_buffer[28]<<1)-(layer_in_buffer[28]<<6)+(layer_in_buffer[28]<<12)+(layer_in_buffer[28]<<14))-(0-(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<12)+(layer_in_buffer[29]<<13))+(0+(layer_in_buffer[30]<<2)-(layer_in_buffer[30]<<4)-(layer_in_buffer[30]<<7)+(layer_in_buffer[30]<<10)+(layer_in_buffer[30]<<12))-(0-(layer_in_buffer[31]<<0)-(layer_in_buffer[31]<<3)-(layer_in_buffer[31]<<5)-(layer_in_buffer[31]<<7)+(layer_in_buffer[31]<<10)+(layer_in_buffer[31]<<13))-(0+(layer_in_buffer[32]<<3)-(layer_in_buffer[32]<<6)+(layer_in_buffer[32]<<11))-(0+(layer_in_buffer[33]<<0)+(layer_in_buffer[33]<<2)-(layer_in_buffer[33]<<4)-(layer_in_buffer[33]<<7)+(layer_in_buffer[33]<<11))+(0-(layer_in_buffer[34]<<3)+(layer_in_buffer[34]<<6)-(layer_in_buffer[34]<<8)+(layer_in_buffer[34]<<10)+(layer_in_buffer[34]<<11)+(layer_in_buffer[34]<<14))-(0+(layer_in_buffer[35]<<1)+(layer_in_buffer[35]<<2)+(layer_in_buffer[35]<<5)+(layer_in_buffer[35]<<7))-(0-(layer_in_buffer[36]<<1)-(layer_in_buffer[36]<<3)-(layer_in_buffer[36]<<5)+(layer_in_buffer[36]<<9)+(layer_in_buffer[36]<<10))-(0+(layer_in_buffer[37]<<0)+(layer_in_buffer[37]<<1)-(layer_in_buffer[37]<<5)+(layer_in_buffer[37]<<7)+(layer_in_buffer[37]<<8)-(layer_in_buffer[37]<<11)+(layer_in_buffer[37]<<14))-(0-(layer_in_buffer[38]<<0)+(layer_in_buffer[38]<<10)+(layer_in_buffer[38]<<11))-(0-(layer_in_buffer[39]<<0)-(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<5)+(layer_in_buffer[39]<<11))+(0+(layer_in_buffer[40]<<1)+(layer_in_buffer[40]<<3)-(layer_in_buffer[40]<<5)-(layer_in_buffer[40]<<8)+(layer_in_buffer[40]<<12))+(0+(layer_in_buffer[41]<<0)+(layer_in_buffer[41]<<5)+(layer_in_buffer[41]<<8)+(layer_in_buffer[41]<<9)+(layer_in_buffer[41]<<12))-(0-(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<3)-(layer_in_buffer[42]<<6)+(layer_in_buffer[42]<<10)+(layer_in_buffer[42]<<12))+(0-(layer_in_buffer[43]<<0)-(layer_in_buffer[43]<<2)+(layer_in_buffer[43]<<5)+(layer_in_buffer[43]<<11))-(0+(layer_in_buffer[44]<<0)+(layer_in_buffer[44]<<2)+(layer_in_buffer[44]<<5)-(layer_in_buffer[44]<<9)-(layer_in_buffer[44]<<11)+(layer_in_buffer[44]<<14))-(0+(layer_in_buffer[45]<<5)+(layer_in_buffer[45]<<6)+(layer_in_buffer[45]<<9)+(layer_in_buffer[45]<<11))+(0+(layer_in_buffer[46]<<1)+(layer_in_buffer[46]<<3)-(layer_in_buffer[46]<<5)-(layer_in_buffer[46]<<8)+(layer_in_buffer[46]<<12))+(0-(layer_in_buffer[47]<<0)-(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<6)-(layer_in_buffer[47]<<8)+(layer_in_buffer[47]<<11)+(layer_in_buffer[47]<<13))-(0+(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<1)+(layer_in_buffer[48]<<4)+(layer_in_buffer[48]<<6))-(0+(layer_in_buffer[49]<<1)-(layer_in_buffer[49]<<3)-(layer_in_buffer[49]<<5)+(layer_in_buffer[49]<<8)+(layer_in_buffer[49]<<11)+(layer_in_buffer[49]<<13))+(0-(layer_in_buffer[50]<<0)+(layer_in_buffer[50]<<3)-(layer_in_buffer[50]<<5)+(layer_in_buffer[50]<<8)+(layer_in_buffer[50]<<9)+(layer_in_buffer[50]<<12)+(layer_in_buffer[50]<<13))-(0+(layer_in_buffer[51]<<0)-(layer_in_buffer[51]<<7)-(layer_in_buffer[51]<<9)+(layer_in_buffer[51]<<13))-(0+(layer_in_buffer[52]<<0)+(layer_in_buffer[52]<<1)-(layer_in_buffer[52]<<4)+(layer_in_buffer[52]<<8)+(layer_in_buffer[52]<<11)+(layer_in_buffer[52]<<14))+(0+(layer_in_buffer[53]<<1)+(layer_in_buffer[53]<<4)+(layer_in_buffer[53]<<6)+(layer_in_buffer[53]<<10)+(layer_in_buffer[53]<<11))-(0+(layer_in_buffer[54]<<0)-(layer_in_buffer[54]<<3)+(layer_in_buffer[54]<<10)+(layer_in_buffer[54]<<12)+(layer_in_buffer[54]<<14))+(0+(layer_in_buffer[55]<<2)+(layer_in_buffer[55]<<4)+(layer_in_buffer[55]<<8)+(layer_in_buffer[55]<<11))+(0+(layer_in_buffer[56]<<0)+(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<3)-(layer_in_buffer[56]<<6)-(layer_in_buffer[56]<<8)+(layer_in_buffer[56]<<13))+(0+(layer_in_buffer[57]<<1)+(layer_in_buffer[57]<<2)+(layer_in_buffer[57]<<5)+(layer_in_buffer[57]<<7))+(0-(layer_in_buffer[58]<<0)+(layer_in_buffer[58]<<4)+(layer_in_buffer[58]<<5)+(layer_in_buffer[58]<<8)+(layer_in_buffer[58]<<12))+(0+(layer_in_buffer[59]<<0)+(layer_in_buffer[59]<<2)+(layer_in_buffer[59]<<3)+(layer_in_buffer[59]<<7)+(layer_in_buffer[59]<<9)+(layer_in_buffer[59]<<10)+(layer_in_buffer[59]<<15))-(0+(layer_in_buffer[60]<<0)-(layer_in_buffer[60]<<2)+(layer_in_buffer[60]<<5)+(layer_in_buffer[60]<<6)-(layer_in_buffer[60]<<9)+(layer_in_buffer[60]<<12)+(layer_in_buffer[60]<<13))-(0+(layer_in_buffer[61]<<0)+(layer_in_buffer[61]<<2)-(layer_in_buffer[61]<<5)-(layer_in_buffer[61]<<9)+(layer_in_buffer[61]<<13)+(layer_in_buffer[61]<<15))+(0-(layer_in_buffer[62]<<2)-(layer_in_buffer[62]<<4)+(layer_in_buffer[62]<<9)+(layer_in_buffer[62]<<11)+(layer_in_buffer[62]<<14))-(0+(layer_in_buffer[63]<<1)+(layer_in_buffer[63]<<3)+(layer_in_buffer[63]<<7)+(layer_in_buffer[63]<<10));
wire [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0-(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<4)-(layer_in_buffer[0]<<7)-(layer_in_buffer[0]<<11)+(layer_in_buffer[0]<<14))-(0+(layer_in_buffer[1]<<7)+(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<11)+(layer_in_buffer[1]<<13))+(0+(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<9))-(0+(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<3)+(layer_in_buffer[3]<<5)+(layer_in_buffer[3]<<9)+(layer_in_buffer[3]<<10))-(0+(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<1)-(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<9)+(layer_in_buffer[4]<<10))-(0-(layer_in_buffer[5]<<2)-(layer_in_buffer[5]<<5)+(layer_in_buffer[5]<<8)+(layer_in_buffer[5]<<12))-(0+(layer_in_buffer[6]<<6)+(layer_in_buffer[6]<<7)+(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<12))-(0+(layer_in_buffer[7]<<7)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<11)+(layer_in_buffer[7]<<13))+(0+(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<5)+(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<9)+(layer_in_buffer[8]<<12))+(0-(layer_in_buffer[9]<<1)+(layer_in_buffer[9]<<6)+(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<9))-(0+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<12)+(layer_in_buffer[10]<<13))-(0-(layer_in_buffer[11]<<1)+(layer_in_buffer[11]<<6)+(layer_in_buffer[11]<<7)-(layer_in_buffer[11]<<10)+(layer_in_buffer[11]<<12)+(layer_in_buffer[11]<<13))+(0+(layer_in_buffer[12]<<0)+(layer_in_buffer[12]<<3)+(layer_in_buffer[12]<<5)+(layer_in_buffer[12]<<9)+(layer_in_buffer[12]<<10))-(0-(layer_in_buffer[13]<<0)-(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<5)+(layer_in_buffer[13]<<11))-(0+(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<4)-(layer_in_buffer[14]<<6)+(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<13))+(0-(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<10)+(layer_in_buffer[15]<<11))-(0+(layer_in_buffer[16]<<0)+(layer_in_buffer[16]<<5)+(layer_in_buffer[16]<<8)+(layer_in_buffer[16]<<9)+(layer_in_buffer[16]<<12))+(0-(layer_in_buffer[17]<<0)+(layer_in_buffer[17]<<5)+(layer_in_buffer[17]<<7)+(layer_in_buffer[17]<<8))+(0+(layer_in_buffer[18]<<5)+(layer_in_buffer[18]<<6)+(layer_in_buffer[18]<<9)+(layer_in_buffer[18]<<11))+(0+(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<6)+(layer_in_buffer[19]<<9)+(layer_in_buffer[19]<<11))-(0-(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<5)+(layer_in_buffer[20]<<6)-(layer_in_buffer[20]<<9)+(layer_in_buffer[20]<<11)+(layer_in_buffer[20]<<12))+(0+(layer_in_buffer[21]<<0)-(layer_in_buffer[21]<<3)-(layer_in_buffer[21]<<5)-(layer_in_buffer[21]<<7)+(layer_in_buffer[21]<<10)+(layer_in_buffer[21]<<11))+(0-(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<8))+(0+(layer_in_buffer[23]<<4)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<10)+(layer_in_buffer[23]<<13))+(0+(layer_in_buffer[24]<<0)+(layer_in_buffer[24]<<2)+(layer_in_buffer[24]<<6)+(layer_in_buffer[24]<<9))+(0+(layer_in_buffer[25]<<2)-(layer_in_buffer[25]<<5)+(layer_in_buffer[25]<<10))+(0-(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<2)-(layer_in_buffer[26]<<4)-(layer_in_buffer[26]<<6)+(layer_in_buffer[26]<<11)+(layer_in_buffer[26]<<12))-(0-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<7)+(layer_in_buffer[27]<<9)+(layer_in_buffer[27]<<10))-(0-(layer_in_buffer[28]<<1)-(layer_in_buffer[28]<<3)-(layer_in_buffer[28]<<5)+(layer_in_buffer[28]<<9)+(layer_in_buffer[28]<<10))+(0-(layer_in_buffer[29]<<0)+(layer_in_buffer[29]<<5)+(layer_in_buffer[29]<<7)+(layer_in_buffer[29]<<8))+(0-(layer_in_buffer[30]<<0)-(layer_in_buffer[30]<<3)+(layer_in_buffer[30]<<6)+(layer_in_buffer[30]<<10))+(0+(layer_in_buffer[31]<<0)+(layer_in_buffer[31]<<1)-(layer_in_buffer[31]<<5)+(layer_in_buffer[31]<<12))+(0+(layer_in_buffer[32]<<1)-(layer_in_buffer[32]<<3)-(layer_in_buffer[32]<<6)+(layer_in_buffer[32]<<9)+(layer_in_buffer[32]<<11))+(0+(layer_in_buffer[33]<<1)+(layer_in_buffer[33]<<2)+(layer_in_buffer[33]<<5)+(layer_in_buffer[33]<<7))-(0+(layer_in_buffer[34]<<2)+(layer_in_buffer[34]<<3)-(layer_in_buffer[34]<<6)-(layer_in_buffer[34]<<8)-(layer_in_buffer[34]<<10)+(layer_in_buffer[34]<<12)+(layer_in_buffer[34]<<13))+(0+(layer_in_buffer[35]<<1)+(layer_in_buffer[35]<<3)+(layer_in_buffer[35]<<7)+(layer_in_buffer[35]<<10))-(0-(layer_in_buffer[36]<<1)+(layer_in_buffer[36]<<6)+(layer_in_buffer[36]<<8)+(layer_in_buffer[36]<<9))-(0-(layer_in_buffer[37]<<0)+(layer_in_buffer[37]<<5)+(layer_in_buffer[37]<<7)+(layer_in_buffer[37]<<8))-(0-(layer_in_buffer[38]<<0)+(layer_in_buffer[38]<<2)+(layer_in_buffer[38]<<3)+(layer_in_buffer[38]<<6)+(layer_in_buffer[38]<<8)+(layer_in_buffer[38]<<10)+(layer_in_buffer[38]<<11))+(0+(layer_in_buffer[39]<<0)+(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<3)+(layer_in_buffer[39]<<9)+(layer_in_buffer[39]<<11))+(0+(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<3)+(layer_in_buffer[40]<<8))-(0+(layer_in_buffer[41]<<2)+(layer_in_buffer[41]<<3)+(layer_in_buffer[41]<<6)+(layer_in_buffer[41]<<8))+(0+(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<2)-(layer_in_buffer[42]<<4)-(layer_in_buffer[42]<<7)+(layer_in_buffer[42]<<11))-(0+(layer_in_buffer[43]<<0)+(layer_in_buffer[43]<<3)+(layer_in_buffer[43]<<9)-(layer_in_buffer[43]<<11)+(layer_in_buffer[43]<<14))+(0+(layer_in_buffer[44]<<0)+(layer_in_buffer[44]<<3)+(layer_in_buffer[44]<<5)+(layer_in_buffer[44]<<9)+(layer_in_buffer[44]<<10))-(0+(layer_in_buffer[45]<<0)+(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<3)+(layer_in_buffer[45]<<9)+(layer_in_buffer[45]<<11))+(0+(layer_in_buffer[46]<<0)+(layer_in_buffer[46]<<3)+(layer_in_buffer[46]<<7)+(layer_in_buffer[46]<<12))+(0+(layer_in_buffer[47]<<2)+(layer_in_buffer[47]<<4)+(layer_in_buffer[47]<<5)+(layer_in_buffer[47]<<11)+(layer_in_buffer[47]<<13))+(0-(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<2)+(layer_in_buffer[48]<<3)+(layer_in_buffer[48]<<6)+(layer_in_buffer[48]<<8)+(layer_in_buffer[48]<<10)+(layer_in_buffer[48]<<11))-(0+(layer_in_buffer[49]<<1)-(layer_in_buffer[49]<<4)-(layer_in_buffer[49]<<6)-(layer_in_buffer[49]<<8)+(layer_in_buffer[49]<<11)+(layer_in_buffer[49]<<12))-(0-(layer_in_buffer[50]<<0)+(layer_in_buffer[50]<<2)+(layer_in_buffer[50]<<3)+(layer_in_buffer[50]<<6)+(layer_in_buffer[50]<<8)+(layer_in_buffer[50]<<10)+(layer_in_buffer[50]<<11))+(0-(layer_in_buffer[51]<<1)+(layer_in_buffer[51]<<4)+(layer_in_buffer[51]<<8)+(layer_in_buffer[51]<<12)+(layer_in_buffer[51]<<14))+(0+(layer_in_buffer[52]<<1)+(layer_in_buffer[52]<<3)+(layer_in_buffer[52]<<7)+(layer_in_buffer[52]<<10))+(0-(layer_in_buffer[53]<<1)-(layer_in_buffer[53]<<4)+(layer_in_buffer[53]<<7)+(layer_in_buffer[53]<<11))+(0+(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<6)-(layer_in_buffer[54]<<9)+(layer_in_buffer[54]<<12))-(0+(layer_in_buffer[55]<<0)+(layer_in_buffer[55]<<1)+(layer_in_buffer[55]<<6)+(layer_in_buffer[55]<<9)+(layer_in_buffer[55]<<11)+(layer_in_buffer[55]<<12))+(0-(layer_in_buffer[56]<<2)+(layer_in_buffer[56]<<7)+(layer_in_buffer[56]<<9)+(layer_in_buffer[56]<<10))-(0-(layer_in_buffer[57]<<0)-(layer_in_buffer[57]<<2)-(layer_in_buffer[57]<<4)+(layer_in_buffer[57]<<8)+(layer_in_buffer[57]<<9))-(0+(layer_in_buffer[58]<<0)+(layer_in_buffer[58]<<1)+(layer_in_buffer[58]<<4)+(layer_in_buffer[58]<<8)+(layer_in_buffer[58]<<10)+(layer_in_buffer[58]<<12))-(0+(layer_in_buffer[59]<<2)+(layer_in_buffer[59]<<4)-(layer_in_buffer[59]<<6)-(layer_in_buffer[59]<<9)+(layer_in_buffer[59]<<13))+(0-(layer_in_buffer[60]<<1)+(layer_in_buffer[60]<<6)+(layer_in_buffer[60]<<8)+(layer_in_buffer[60]<<9))-(0+(layer_in_buffer[61]<<1)+(layer_in_buffer[61]<<3)+(layer_in_buffer[61]<<7)+(layer_in_buffer[61]<<10))+(0-(layer_in_buffer[62]<<1)-(layer_in_buffer[62]<<3)-(layer_in_buffer[62]<<5)+(layer_in_buffer[62]<<9)+(layer_in_buffer[62]<<10))-(0+(layer_in_buffer[63]<<3)+(layer_in_buffer[63]<<4)+(layer_in_buffer[63]<<7)+(layer_in_buffer[63]<<9));
wire [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0+(0+(layer_in_buffer[0]<<0)-(layer_in_buffer[0]<<2)+(layer_in_buffer[0]<<6)-(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<12))-(0-(layer_in_buffer[1]<<0)-(layer_in_buffer[1]<<2)-(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<8)-(layer_in_buffer[1]<<10)+(layer_in_buffer[1]<<13))-(0-(layer_in_buffer[2]<<0)-(layer_in_buffer[2]<<2)+(layer_in_buffer[2]<<5)+(layer_in_buffer[2]<<11))-(0-(layer_in_buffer[3]<<0)+(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<3)+(layer_in_buffer[3]<<6)+(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<11))+(0+(layer_in_buffer[4]<<1)+(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<8)+(layer_in_buffer[4]<<10)+(layer_in_buffer[4]<<11))-(0+(layer_in_buffer[5]<<0)+(layer_in_buffer[5]<<2)-(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<8)+(layer_in_buffer[5]<<12)+(layer_in_buffer[5]<<13))+(0+(layer_in_buffer[6]<<1)-(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<7)-(layer_in_buffer[6]<<9)+(layer_in_buffer[6]<<13))+(0+(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<1)-(layer_in_buffer[7]<<4)-(layer_in_buffer[7]<<6)-(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<10)+(layer_in_buffer[7]<<11))-(0+(layer_in_buffer[8]<<1)-(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<12)+(layer_in_buffer[8]<<14))-(0-(layer_in_buffer[9]<<1)-(layer_in_buffer[9]<<3)+(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<10)+(layer_in_buffer[9]<<13))+(0+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<8)+(layer_in_buffer[10]<<12))-(0+(layer_in_buffer[11]<<0)-(layer_in_buffer[11]<<3)+(layer_in_buffer[11]<<6)+(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<12)+(layer_in_buffer[11]<<15))-(0-(layer_in_buffer[12]<<0)-(layer_in_buffer[12]<<2)-(layer_in_buffer[12]<<4)-(layer_in_buffer[12]<<6)+(layer_in_buffer[12]<<11)+(layer_in_buffer[12]<<12))+(0+(layer_in_buffer[13]<<0)+(layer_in_buffer[13]<<2)+(layer_in_buffer[13]<<6)+(layer_in_buffer[13]<<9))+(0-(layer_in_buffer[14]<<0)-(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<9)+(layer_in_buffer[14]<<10)+(layer_in_buffer[14]<<13))-(0-(layer_in_buffer[15]<<0)-(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<10))-(0-(layer_in_buffer[16]<<2)-(layer_in_buffer[16]<<4)+(layer_in_buffer[16]<<7)+(layer_in_buffer[16]<<13))+(0-(layer_in_buffer[17]<<0)-(layer_in_buffer[17]<<2)-(layer_in_buffer[17]<<5)+(layer_in_buffer[17]<<8)-(layer_in_buffer[17]<<10)+(layer_in_buffer[17]<<13))-(0+(layer_in_buffer[18]<<1)+(layer_in_buffer[18]<<3)+(layer_in_buffer[18]<<6)+(layer_in_buffer[18]<<8)+(layer_in_buffer[18]<<11)+(layer_in_buffer[18]<<12))-(0-(layer_in_buffer[19]<<2)-(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<8)+(layer_in_buffer[19]<<12))-(0+(layer_in_buffer[20]<<0)+(layer_in_buffer[20]<<2)+(layer_in_buffer[20]<<6)+(layer_in_buffer[20]<<9))+(0-(layer_in_buffer[21]<<3)+(layer_in_buffer[21]<<8)+(layer_in_buffer[21]<<10)+(layer_in_buffer[21]<<11))-(0+(layer_in_buffer[22]<<3)+(layer_in_buffer[22]<<5)+(layer_in_buffer[22]<<9)+(layer_in_buffer[22]<<12))+(0+(layer_in_buffer[23]<<0)+(layer_in_buffer[23]<<6)+(layer_in_buffer[23]<<7)+(layer_in_buffer[23]<<11))+(0-(layer_in_buffer[24]<<1)+(layer_in_buffer[24]<<6)+(layer_in_buffer[24]<<8)+(layer_in_buffer[24]<<9))-(0+(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<1)+(layer_in_buffer[25]<<4)+(layer_in_buffer[25]<<5)+(layer_in_buffer[25]<<10)+(layer_in_buffer[25]<<12)+(layer_in_buffer[25]<<13))+(0+(layer_in_buffer[26]<<1)+(layer_in_buffer[26]<<3)-(layer_in_buffer[26]<<5)-(layer_in_buffer[26]<<8)+(layer_in_buffer[26]<<12))+(0-(layer_in_buffer[28]<<3)+(layer_in_buffer[28]<<8)+(layer_in_buffer[28]<<10)+(layer_in_buffer[28]<<11))-(0-(layer_in_buffer[29]<<0)+(layer_in_buffer[29]<<3)-(layer_in_buffer[29]<<5)+(layer_in_buffer[29]<<7)+(layer_in_buffer[29]<<8)+(layer_in_buffer[29]<<11))+(0+(layer_in_buffer[30]<<5)+(layer_in_buffer[30]<<6)+(layer_in_buffer[30]<<9)+(layer_in_buffer[30]<<11))+(0+(layer_in_buffer[31]<<1)+(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<6)+(layer_in_buffer[31]<<10)+(layer_in_buffer[31]<<11))+(0-(layer_in_buffer[32]<<0)-(layer_in_buffer[32]<<2)+(layer_in_buffer[32]<<5)+(layer_in_buffer[32]<<11))+(0+(layer_in_buffer[33]<<0)+(layer_in_buffer[33]<<1)-(layer_in_buffer[33]<<4)-(layer_in_buffer[33]<<6)-(layer_in_buffer[33]<<8)+(layer_in_buffer[33]<<10)+(layer_in_buffer[33]<<11))+(0+(layer_in_buffer[34]<<0)+(layer_in_buffer[34]<<4)+(layer_in_buffer[34]<<6)+(layer_in_buffer[34]<<11)+(layer_in_buffer[34]<<12))+(0-(layer_in_buffer[35]<<1)+(layer_in_buffer[35]<<6)+(layer_in_buffer[35]<<8)+(layer_in_buffer[35]<<9))+(0-(layer_in_buffer[36]<<1)-(layer_in_buffer[36]<<3)-(layer_in_buffer[36]<<5)+(layer_in_buffer[36]<<9)+(layer_in_buffer[36]<<10))+(0-(layer_in_buffer[37]<<1)+(layer_in_buffer[37]<<4)+(layer_in_buffer[37]<<5)+(layer_in_buffer[37]<<8)-(layer_in_buffer[37]<<10)+(layer_in_buffer[37]<<13))+(0+(layer_in_buffer[38]<<1)-(layer_in_buffer[38]<<4)+(layer_in_buffer[38]<<9))+(0+(layer_in_buffer[39]<<0)+(layer_in_buffer[39]<<2)+(layer_in_buffer[39]<<6)+(layer_in_buffer[39]<<9))-(0+(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<4)+(layer_in_buffer[40]<<7)+(layer_in_buffer[40]<<9)+(layer_in_buffer[40]<<11)+(layer_in_buffer[40]<<15))+(0+(layer_in_buffer[41]<<0)+(layer_in_buffer[41]<<1)-(layer_in_buffer[41]<<7)+(layer_in_buffer[41]<<9)+(layer_in_buffer[41]<<10))-(0-(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<2)+(layer_in_buffer[42]<<3)-(layer_in_buffer[42]<<7)+(layer_in_buffer[42]<<10)+(layer_in_buffer[42]<<11)+(layer_in_buffer[42]<<14))+(0-(layer_in_buffer[43]<<0)+(layer_in_buffer[43]<<4)-(layer_in_buffer[43]<<6)-(layer_in_buffer[43]<<8)+(layer_in_buffer[43]<<11))+(0-(layer_in_buffer[44]<<1)+(layer_in_buffer[44]<<5)-(layer_in_buffer[44]<<7)-(layer_in_buffer[44]<<9)+(layer_in_buffer[44]<<12))-(0+(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6)+(layer_in_buffer[45]<<8)+(layer_in_buffer[45]<<13)+(layer_in_buffer[45]<<14))-(0+(layer_in_buffer[46]<<2)+(layer_in_buffer[46]<<3)+(layer_in_buffer[46]<<6)+(layer_in_buffer[46]<<8))-(0+(layer_in_buffer[47]<<1)-(layer_in_buffer[47]<<3)+(layer_in_buffer[47]<<6)+(layer_in_buffer[47]<<8)+(layer_in_buffer[47]<<9)+(layer_in_buffer[47]<<12)+(layer_in_buffer[47]<<13))+(0+(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<2)+(layer_in_buffer[48]<<6)+(layer_in_buffer[48]<<9))+(0+(layer_in_buffer[49]<<1)+(layer_in_buffer[49]<<2)+(layer_in_buffer[49]<<7)+(layer_in_buffer[49]<<10)+(layer_in_buffer[49]<<12)+(layer_in_buffer[49]<<13))-(0-(layer_in_buffer[50]<<0)+(layer_in_buffer[50]<<4)-(layer_in_buffer[50]<<6)+(layer_in_buffer[50]<<9)-(layer_in_buffer[50]<<11)+(layer_in_buffer[50]<<13)+(layer_in_buffer[50]<<14))+(0+(layer_in_buffer[51]<<3)+(layer_in_buffer[51]<<7)-(layer_in_buffer[51]<<10)+(layer_in_buffer[51]<<13))+(0+(layer_in_buffer[52]<<0)+(layer_in_buffer[52]<<6)+(layer_in_buffer[52]<<7)+(layer_in_buffer[52]<<11))+(0-(layer_in_buffer[53]<<1)-(layer_in_buffer[53]<<3)-(layer_in_buffer[53]<<5)+(layer_in_buffer[53]<<9)+(layer_in_buffer[53]<<10))+(0+(layer_in_buffer[54]<<1)+(layer_in_buffer[54]<<4)+(layer_in_buffer[54]<<6)+(layer_in_buffer[54]<<10)+(layer_in_buffer[54]<<11))+(0+(layer_in_buffer[55]<<1)-(layer_in_buffer[55]<<4)+(layer_in_buffer[55]<<9))-(0-(layer_in_buffer[56]<<1)+(layer_in_buffer[56]<<6)-(layer_in_buffer[56]<<9)-(layer_in_buffer[56]<<11)+(layer_in_buffer[56]<<13)+(layer_in_buffer[56]<<14))+(0+(layer_in_buffer[57]<<3)+(layer_in_buffer[57]<<7)-(layer_in_buffer[57]<<10)+(layer_in_buffer[57]<<13))+(0+(layer_in_buffer[58]<<2)+(layer_in_buffer[58]<<8)+(layer_in_buffer[58]<<9)+(layer_in_buffer[58]<<13))-(0-(layer_in_buffer[59]<<0)+(layer_in_buffer[59]<<3)+(layer_in_buffer[59]<<5)-(layer_in_buffer[59]<<9)+(layer_in_buffer[59]<<13))-(0-(layer_in_buffer[60]<<3)+(layer_in_buffer[60]<<8)+(layer_in_buffer[60]<<10)+(layer_in_buffer[60]<<11))-(0+(layer_in_buffer[61]<<0)+(layer_in_buffer[61]<<2)-(layer_in_buffer[61]<<4)-(layer_in_buffer[61]<<6)+(layer_in_buffer[61]<<9)+(layer_in_buffer[61]<<10)+(layer_in_buffer[61]<<14))-(0+(layer_in_buffer[62]<<2)+(layer_in_buffer[62]<<5)+(layer_in_buffer[62]<<6)+(layer_in_buffer[62]<<15))+(0-(layer_in_buffer[63]<<1)+(layer_in_buffer[63]<<6)+(layer_in_buffer[63]<<8)+(layer_in_buffer[63]<<9));
wire [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0+(0+(layer_in_buffer[0]<<1)+(layer_in_buffer[0]<<4)+(layer_in_buffer[0]<<6)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<11))+(0+(layer_in_buffer[1]<<1)+(layer_in_buffer[1]<<5)-(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<11))+(0+(layer_in_buffer[2]<<0)+(layer_in_buffer[2]<<1)+(layer_in_buffer[2]<<4)+(layer_in_buffer[2]<<8)+(layer_in_buffer[2]<<10)+(layer_in_buffer[2]<<12))-(0+(layer_in_buffer[3]<<1)+(layer_in_buffer[3]<<3)+(layer_in_buffer[3]<<5)-(layer_in_buffer[3]<<7)+(layer_in_buffer[3]<<10)+(layer_in_buffer[3]<<13))+(0+(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<6)+(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<11))+(0+(layer_in_buffer[5]<<0)-(layer_in_buffer[5]<<2)+(layer_in_buffer[5]<<4)+(layer_in_buffer[5]<<5)+(layer_in_buffer[5]<<8)+(layer_in_buffer[5]<<11)+(layer_in_buffer[5]<<13))+(0-(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<3)+(layer_in_buffer[6]<<4)+(layer_in_buffer[6]<<7)-(layer_in_buffer[6]<<9)+(layer_in_buffer[6]<<12))-(0+(layer_in_buffer[7]<<1)+(layer_in_buffer[7]<<3)-(layer_in_buffer[7]<<6)+(layer_in_buffer[7]<<8)+(layer_in_buffer[7]<<9)+(layer_in_buffer[7]<<14))-(0+(layer_in_buffer[8]<<4)+(layer_in_buffer[8]<<5)+(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<10))+(0+(layer_in_buffer[9]<<1)-(layer_in_buffer[9]<<3)-(layer_in_buffer[9]<<6)+(layer_in_buffer[9]<<9)+(layer_in_buffer[9]<<11))+(0+(layer_in_buffer[10]<<1)+(layer_in_buffer[10]<<2)+(layer_in_buffer[10]<<5)+(layer_in_buffer[10]<<7))-(0-(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<3)+(layer_in_buffer[11]<<4)+(layer_in_buffer[11]<<7)-(layer_in_buffer[11]<<9)+(layer_in_buffer[11]<<12))+(0-(layer_in_buffer[12]<<3)+(layer_in_buffer[12]<<8)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<11))+(0-(layer_in_buffer[13]<<3)+(layer_in_buffer[13]<<8)+(layer_in_buffer[13]<<10)+(layer_in_buffer[13]<<11))+(0+(layer_in_buffer[14]<<0)+(layer_in_buffer[14]<<2)-(layer_in_buffer[14]<<5)-(layer_in_buffer[14]<<8)+(layer_in_buffer[14]<<10)+(layer_in_buffer[14]<<11)+(layer_in_buffer[14]<<14))+(0-(layer_in_buffer[15]<<0)+(layer_in_buffer[15]<<4)-(layer_in_buffer[15]<<6)-(layer_in_buffer[15]<<8)+(layer_in_buffer[15]<<11))+(0+(layer_in_buffer[16]<<0)+(layer_in_buffer[16]<<1)-(layer_in_buffer[16]<<5)+(layer_in_buffer[16]<<12))-(0+(layer_in_buffer[17]<<0)+(layer_in_buffer[17]<<1)+(layer_in_buffer[17]<<4)+(layer_in_buffer[17]<<7)-(layer_in_buffer[17]<<9)+(layer_in_buffer[17]<<14))+(0+(layer_in_buffer[18]<<1)+(layer_in_buffer[18]<<5)-(layer_in_buffer[18]<<8)+(layer_in_buffer[18]<<11))+(0-(layer_in_buffer[19]<<1)+(layer_in_buffer[19]<<6)+(layer_in_buffer[19]<<8)+(layer_in_buffer[19]<<9))+(0-(layer_in_buffer[20]<<3)+(layer_in_buffer[20]<<8)+(layer_in_buffer[20]<<10)+(layer_in_buffer[20]<<11))+(0+(layer_in_buffer[21]<<1)+(layer_in_buffer[21]<<5)-(layer_in_buffer[21]<<8)+(layer_in_buffer[21]<<11))+(0+(layer_in_buffer[22]<<0)+(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<6)+(layer_in_buffer[22]<<9))+(0-(layer_in_buffer[23]<<0)-(layer_in_buffer[23]<<4)+(layer_in_buffer[23]<<9)+(layer_in_buffer[23]<<10)+(layer_in_buffer[23]<<13))-(0+(layer_in_buffer[24]<<3)+(layer_in_buffer[24]<<4)+(layer_in_buffer[24]<<7)+(layer_in_buffer[24]<<9))+(0+(layer_in_buffer[25]<<2)+(layer_in_buffer[25]<<4)+(layer_in_buffer[25]<<8)+(layer_in_buffer[25]<<11))-(0-(layer_in_buffer[26]<<0)-(layer_in_buffer[26]<<4)+(layer_in_buffer[26]<<9)+(layer_in_buffer[26]<<10)+(layer_in_buffer[26]<<13))-(0-(layer_in_buffer[27]<<2)+(layer_in_buffer[27]<<6)-(layer_in_buffer[27]<<9)-(layer_in_buffer[27]<<12)+(layer_in_buffer[27]<<15))+(0+(layer_in_buffer[28]<<0)+(layer_in_buffer[28]<<4)-(layer_in_buffer[28]<<7)+(layer_in_buffer[28]<<10))+(0-(layer_in_buffer[29]<<0)+(layer_in_buffer[29]<<3)+(layer_in_buffer[29]<<4)+(layer_in_buffer[29]<<7)-(layer_in_buffer[29]<<9)+(layer_in_buffer[29]<<12))-(0+(layer_in_buffer[30]<<3)-(layer_in_buffer[30]<<5)-(layer_in_buffer[30]<<8)+(layer_in_buffer[30]<<11)+(layer_in_buffer[30]<<13))+(0+(layer_in_buffer[31]<<6)+(layer_in_buffer[31]<<7)+(layer_in_buffer[31]<<10)+(layer_in_buffer[31]<<12))+(0+(layer_in_buffer[32]<<0)+(layer_in_buffer[32]<<6)+(layer_in_buffer[32]<<7)+(layer_in_buffer[32]<<11))+(0+(layer_in_buffer[33]<<0)+(layer_in_buffer[33]<<3)+(layer_in_buffer[33]<<5)+(layer_in_buffer[33]<<9)+(layer_in_buffer[33]<<10))+(0+(layer_in_buffer[34]<<3)+(layer_in_buffer[34]<<5)+(layer_in_buffer[34]<<9)+(layer_in_buffer[34]<<12))-(0-(layer_in_buffer[35]<<0)-(layer_in_buffer[35]<<2)-(layer_in_buffer[35]<<4)+(layer_in_buffer[35]<<8)+(layer_in_buffer[35]<<9))+(0+(layer_in_buffer[36]<<0)+(layer_in_buffer[36]<<1)+(layer_in_buffer[36]<<6)+(layer_in_buffer[36]<<9)+(layer_in_buffer[36]<<11)+(layer_in_buffer[36]<<12))-(0+(layer_in_buffer[37]<<1)+(layer_in_buffer[37]<<4)+(layer_in_buffer[37]<<6)+(layer_in_buffer[37]<<10)+(layer_in_buffer[37]<<11))-(0+(layer_in_buffer[38]<<1)+(layer_in_buffer[38]<<2)+(layer_in_buffer[38]<<5)+(layer_in_buffer[38]<<9)+(layer_in_buffer[38]<<11)+(layer_in_buffer[38]<<13))+(0+(layer_in_buffer[39]<<0)+(layer_in_buffer[39]<<2)-(layer_in_buffer[39]<<4)-(layer_in_buffer[39]<<7)+(layer_in_buffer[39]<<11))-(0+(layer_in_buffer[40]<<0)+(layer_in_buffer[40]<<1)-(layer_in_buffer[40]<<7)+(layer_in_buffer[40]<<9)+(layer_in_buffer[40]<<10))+(0+(layer_in_buffer[41]<<5)+(layer_in_buffer[41]<<6)+(layer_in_buffer[41]<<9)+(layer_in_buffer[41]<<11))-(0-(layer_in_buffer[42]<<3)+(layer_in_buffer[42]<<8)+(layer_in_buffer[42]<<10)+(layer_in_buffer[42]<<11))+(0+(layer_in_buffer[43]<<2)+(layer_in_buffer[43]<<4)-(layer_in_buffer[43]<<6)-(layer_in_buffer[43]<<9)+(layer_in_buffer[43]<<13))+(0+(layer_in_buffer[44]<<2)+(layer_in_buffer[44]<<4)+(layer_in_buffer[44]<<8)+(layer_in_buffer[44]<<11))-(0-(layer_in_buffer[45]<<2)+(layer_in_buffer[45]<<6)-(layer_in_buffer[45]<<8)-(layer_in_buffer[45]<<10)+(layer_in_buffer[45]<<13))+(0-(layer_in_buffer[46]<<0)+(layer_in_buffer[46]<<5)+(layer_in_buffer[46]<<7)+(layer_in_buffer[46]<<8))-(0+(layer_in_buffer[47]<<0)+(layer_in_buffer[47]<<4)+(layer_in_buffer[47]<<7)-(layer_in_buffer[47]<<9)-(layer_in_buffer[47]<<11)+(layer_in_buffer[47]<<13)+(layer_in_buffer[47]<<14))+(0+(layer_in_buffer[48]<<0)+(layer_in_buffer[48]<<4)-(layer_in_buffer[48]<<7)+(layer_in_buffer[48]<<10))+(0-(layer_in_buffer[49]<<4)-(layer_in_buffer[49]<<6)-(layer_in_buffer[49]<<8)+(layer_in_buffer[49]<<12)+(layer_in_buffer[49]<<13))+(0+(layer_in_buffer[50]<<5)-(layer_in_buffer[50]<<8)+(layer_in_buffer[50]<<13))-(0+(layer_in_buffer[51]<<3)+(layer_in_buffer[51]<<7)+(layer_in_buffer[51]<<9)+(layer_in_buffer[51]<<14)+(layer_in_buffer[51]<<15))-(0+(layer_in_buffer[52]<<0)+(layer_in_buffer[52]<<1)-(layer_in_buffer[52]<<5)+(layer_in_buffer[52]<<12))-(0-(layer_in_buffer[53]<<1)+(layer_in_buffer[53]<<6)+(layer_in_buffer[53]<<8)+(layer_in_buffer[53]<<9))-(0-(layer_in_buffer[54]<<2)+(layer_in_buffer[54]<<7)+(layer_in_buffer[54]<<9)+(layer_in_buffer[54]<<10))+(0+(layer_in_buffer[55]<<0)+(layer_in_buffer[55]<<1)-(layer_in_buffer[55]<<7)+(layer_in_buffer[55]<<9)+(layer_in_buffer[55]<<10))-(0+(layer_in_buffer[56]<<1)+(layer_in_buffer[56]<<2)-(layer_in_buffer[56]<<5)-(layer_in_buffer[56]<<7)-(layer_in_buffer[56]<<9)+(layer_in_buffer[56]<<11)+(layer_in_buffer[56]<<12))-(0+(layer_in_buffer[57]<<0)+(layer_in_buffer[57]<<1)+(layer_in_buffer[57]<<4)+(layer_in_buffer[57]<<7)-(layer_in_buffer[57]<<9)+(layer_in_buffer[57]<<14))+(0+(layer_in_buffer[58]<<0)+(layer_in_buffer[58]<<2)-(layer_in_buffer[58]<<4)-(layer_in_buffer[58]<<7)+(layer_in_buffer[58]<<11))-(0+(layer_in_buffer[59]<<2)-(layer_in_buffer[59]<<5)-(layer_in_buffer[59]<<7)-(layer_in_buffer[59]<<9)+(layer_in_buffer[59]<<12)+(layer_in_buffer[59]<<13))+(0-(layer_in_buffer[60]<<1)+(layer_in_buffer[60]<<5)-(layer_in_buffer[60]<<7)-(layer_in_buffer[60]<<9)+(layer_in_buffer[60]<<12))-(0+(layer_in_buffer[61]<<0)+(layer_in_buffer[61]<<2)-(layer_in_buffer[61]<<4)-(layer_in_buffer[61]<<7)+(layer_in_buffer[61]<<11))-(0+(layer_in_buffer[62]<<1)+(layer_in_buffer[62]<<7)+(layer_in_buffer[62]<<8)+(layer_in_buffer[62]<<12))+(0+(layer_in_buffer[63]<<3)+(layer_in_buffer[63]<<4)+(layer_in_buffer[63]<<7)+(layer_in_buffer[63]<<9));
wire [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0-(0+(layer_in_buffer[0]<<1)+(layer_in_buffer[0]<<2)-(layer_in_buffer[0]<<8)+(layer_in_buffer[0]<<10)+(layer_in_buffer[0]<<11))-(0+(layer_in_buffer[1]<<0)+(layer_in_buffer[1]<<5)+(layer_in_buffer[1]<<8)+(layer_in_buffer[1]<<9)+(layer_in_buffer[1]<<12))-(0+(layer_in_buffer[2]<<1)-(layer_in_buffer[2]<<6)+(layer_in_buffer[2]<<12)+(layer_in_buffer[2]<<14))+(0+(layer_in_buffer[3]<<0)-(layer_in_buffer[3]<<2)+(layer_in_buffer[3]<<6)-(layer_in_buffer[3]<<8)+(layer_in_buffer[3]<<12))-(0+(layer_in_buffer[4]<<0)+(layer_in_buffer[4]<<2)-(layer_in_buffer[4]<<4)-(layer_in_buffer[4]<<7)+(layer_in_buffer[4]<<11))+(0+(layer_in_buffer[5]<<2)-(layer_in_buffer[5]<<4)-(layer_in_buffer[5]<<7)+(layer_in_buffer[5]<<10)+(layer_in_buffer[5]<<12))+(0-(layer_in_buffer[6]<<0)+(layer_in_buffer[6]<<5)-(layer_in_buffer[6]<<8)-(layer_in_buffer[6]<<10)+(layer_in_buffer[6]<<12)+(layer_in_buffer[6]<<13))+(0+(layer_in_buffer[7]<<0)+(layer_in_buffer[7]<<1)-(layer_in_buffer[7]<<5)+(layer_in_buffer[7]<<12))-(0-(layer_in_buffer[8]<<0)+(layer_in_buffer[8]<<2)+(layer_in_buffer[8]<<3)+(layer_in_buffer[8]<<6)+(layer_in_buffer[8]<<8)+(layer_in_buffer[8]<<10)+(layer_in_buffer[8]<<11))-(0+(layer_in_buffer[9]<<0)+(layer_in_buffer[9]<<1)-(layer_in_buffer[9]<<8)+(layer_in_buffer[9]<<12)+(layer_in_buffer[9]<<13))+(0+(layer_in_buffer[10]<<0)-(layer_in_buffer[10]<<2)-(layer_in_buffer[10]<<4)+(layer_in_buffer[10]<<7)+(layer_in_buffer[10]<<10)+(layer_in_buffer[10]<<12))-(0-(layer_in_buffer[11]<<0)+(layer_in_buffer[11]<<4)-(layer_in_buffer[11]<<7)-(layer_in_buffer[11]<<10)+(layer_in_buffer[11]<<13))-(0+(layer_in_buffer[12]<<1)+(layer_in_buffer[12]<<2)-(layer_in_buffer[12]<<8)+(layer_in_buffer[12]<<10)+(layer_in_buffer[12]<<11))+(0-(layer_in_buffer[13]<<1)-(layer_in_buffer[13]<<3)-(layer_in_buffer[13]<<5)+(layer_in_buffer[13]<<9)+(layer_in_buffer[13]<<10))-(0-(layer_in_buffer[14]<<1)+(layer_in_buffer[14]<<4)+(layer_in_buffer[14]<<5)+(layer_in_buffer[14]<<8)-(layer_in_buffer[14]<<10)+(layer_in_buffer[14]<<13))+(0+(layer_in_buffer[15]<<2)+(layer_in_buffer[15]<<3)+(layer_in_buffer[15]<<6)+(layer_in_buffer[15]<<8))+(0+(layer_in_buffer[16]<<4)-(layer_in_buffer[16]<<7)+(layer_in_buffer[16]<<12))-(0+(layer_in_buffer[17]<<0)+(layer_in_buffer[17]<<2)+(layer_in_buffer[17]<<5)-(layer_in_buffer[17]<<9)-(layer_in_buffer[17]<<11)+(layer_in_buffer[17]<<14))+(0-(layer_in_buffer[18]<<0)-(layer_in_buffer[18]<<2)+(layer_in_buffer[18]<<5)+(layer_in_buffer[18]<<11))-(0-(layer_in_buffer[19]<<0)-(layer_in_buffer[19]<<2)+(layer_in_buffer[19]<<5)+(layer_in_buffer[19]<<11))+(0+(layer_in_buffer[20]<<1)+(layer_in_buffer[20]<<7)+(layer_in_buffer[20]<<8)+(layer_in_buffer[20]<<12))+(0-(layer_in_buffer[21]<<0)+(layer_in_buffer[21]<<10)+(layer_in_buffer[21]<<11))-(0-(layer_in_buffer[22]<<0)-(layer_in_buffer[22]<<2)+(layer_in_buffer[22]<<7)+(layer_in_buffer[22]<<9)+(layer_in_buffer[22]<<12))-(0+(layer_in_buffer[23]<<1)+(layer_in_buffer[23]<<5)+(layer_in_buffer[23]<<9)-(layer_in_buffer[23]<<11)+(layer_in_buffer[23]<<13)+(layer_in_buffer[23]<<14))-(0+(layer_in_buffer[24]<<0)+(layer_in_buffer[24]<<1)+(layer_in_buffer[24]<<4)+(layer_in_buffer[24]<<6))-(0-(layer_in_buffer[25]<<0)+(layer_in_buffer[25]<<3)+(layer_in_buffer[25]<<5)-(layer_in_buffer[25]<<9)+(layer_in_buffer[25]<<13))+(0-(layer_in_buffer[26]<<1)+(layer_in_buffer[26]<<5)-(layer_in_buffer[26]<<7)-(layer_in_buffer[26]<<9)+(layer_in_buffer[26]<<12))-(0-(layer_in_buffer[27]<<3)-(layer_in_buffer[27]<<5)-(layer_in_buffer[27]<<7)+(layer_in_buffer[27]<<11)+(layer_in_buffer[27]<<12))-(0-(layer_in_buffer[28]<<2)-(layer_in_buffer[28]<<5)+(layer_in_buffer[28]<<8)+(layer_in_buffer[28]<<12))-(0+(layer_in_buffer[29]<<2)+(layer_in_buffer[29]<<3)+(layer_in_buffer[29]<<6)+(layer_in_buffer[29]<<8))+(0+(layer_in_buffer[30]<<0)+(layer_in_buffer[30]<<2)+(layer_in_buffer[30]<<4)-(layer_in_buffer[30]<<6)+(layer_in_buffer[30]<<9)+(layer_in_buffer[30]<<12))-(0+(layer_in_buffer[31]<<0)+(layer_in_buffer[31]<<1)+(layer_in_buffer[31]<<4)+(layer_in_buffer[31]<<6))+(0+(layer_in_buffer[32]<<0)+(layer_in_buffer[32]<<6)+(layer_in_buffer[32]<<7)+(layer_in_buffer[32]<<11))+(0+(layer_in_buffer[33]<<0)-(layer_in_buffer[33]<<2)+(layer_in_buffer[33]<<6)-(layer_in_buffer[33]<<8)+(layer_in_buffer[33]<<12))-(0+(layer_in_buffer[34]<<1)+(layer_in_buffer[34]<<3)-(layer_in_buffer[34]<<5)+(layer_in_buffer[34]<<9)+(layer_in_buffer[34]<<13)+(layer_in_buffer[34]<<14))+(0+(layer_in_buffer[35]<<0)+(layer_in_buffer[35]<<1)+(layer_in_buffer[35]<<4)+(layer_in_buffer[35]<<6))+(0-(layer_in_buffer[36]<<0)+(layer_in_buffer[36]<<10)+(layer_in_buffer[36]<<11))+(0+(layer_in_buffer[37]<<0)-(layer_in_buffer[37]<<2)-(layer_in_buffer[37]<<5)+(layer_in_buffer[37]<<8)+(layer_in_buffer[37]<<10))+(0+(layer_in_buffer[38]<<0)+(layer_in_buffer[38]<<2)-(layer_in_buffer[38]<<8)+(layer_in_buffer[38]<<11)+(layer_in_buffer[38]<<12))-(0-(layer_in_buffer[39]<<0)-(layer_in_buffer[39]<<2)-(layer_in_buffer[39]<<4)+(layer_in_buffer[39]<<8)+(layer_in_buffer[39]<<9))+(0+(layer_in_buffer[40]<<0)-(layer_in_buffer[40]<<3)-(layer_in_buffer[40]<<6)-(layer_in_buffer[40]<<9)+(layer_in_buffer[40]<<11)+(layer_in_buffer[40]<<12))-(0+(layer_in_buffer[41]<<1)-(layer_in_buffer[41]<<3)-(layer_in_buffer[41]<<6)+(layer_in_buffer[41]<<9)+(layer_in_buffer[41]<<11))-(0-(layer_in_buffer[42]<<0)+(layer_in_buffer[42]<<3)+(layer_in_buffer[42]<<4)+(layer_in_buffer[42]<<7)-(layer_in_buffer[42]<<9)+(layer_in_buffer[42]<<12))+(0-(layer_in_buffer[43]<<1)+(layer_in_buffer[43]<<6)+(layer_in_buffer[43]<<8)+(layer_in_buffer[43]<<9))-(0-(layer_in_buffer[44]<<0)+(layer_in_buffer[44]<<5)-(layer_in_buffer[44]<<8)-(layer_in_buffer[44]<<10)+(layer_in_buffer[44]<<12)+(layer_in_buffer[44]<<13))-(0-(layer_in_buffer[45]<<5)+(layer_in_buffer[45]<<10)+(layer_in_buffer[45]<<12)+(layer_in_buffer[45]<<13))+(0+(layer_in_buffer[46]<<2)+(layer_in_buffer[46]<<4)+(layer_in_buffer[46]<<8)+(layer_in_buffer[46]<<11))-(0-(layer_in_buffer[47]<<1)+(layer_in_buffer[47]<<4)+(layer_in_buffer[47]<<6)-(layer_in_buffer[47]<<10)+(layer_in_buffer[47]<<14))+(0+(layer_in_buffer[48]<<5)+(layer_in_buffer[48]<<6)+(layer_in_buffer[48]<<9)+(layer_in_buffer[48]<<11))-(0+(layer_in_buffer[49]<<0)+(layer_in_buffer[49]<<2)-(layer_in_buffer[49]<<5)+(layer_in_buffer[49]<<7)+(layer_in_buffer[49]<<8)+(layer_in_buffer[49]<<13))-(0-(layer_in_buffer[50]<<0)+(layer_in_buffer[50]<<5)+(layer_in_buffer[50]<<6)-(layer_in_buffer[50]<<9)+(layer_in_buffer[50]<<11)+(layer_in_buffer[50]<<12))+(0+(layer_in_buffer[51]<<0)+(layer_in_buffer[51]<<1)-(layer_in_buffer[51]<<4)-(layer_in_buffer[51]<<6)-(layer_in_buffer[51]<<8)+(layer_in_buffer[51]<<10)+(layer_in_buffer[51]<<11))-(0+(layer_in_buffer[52]<<3)-(layer_in_buffer[52]<<6)+(layer_in_buffer[52]<<11))+(0-(layer_in_buffer[53]<<3)+(layer_in_buffer[53]<<8)+(layer_in_buffer[53]<<10)+(layer_in_buffer[53]<<11))-(0+(layer_in_buffer[54]<<1)+(layer_in_buffer[54]<<4)+(layer_in_buffer[54]<<8)+(layer_in_buffer[54]<<13))+(0+(layer_in_buffer[55]<<1)+(layer_in_buffer[55]<<4)+(layer_in_buffer[55]<<6)+(layer_in_buffer[55]<<10)+(layer_in_buffer[55]<<11))-(0-(layer_in_buffer[56]<<0)+(layer_in_buffer[56]<<4)-(layer_in_buffer[56]<<7)-(layer_in_buffer[56]<<10)+(layer_in_buffer[56]<<13))+(0-(layer_in_buffer[57]<<0)+(layer_in_buffer[57]<<5)+(layer_in_buffer[57]<<7)+(layer_in_buffer[57]<<8))-(0+(layer_in_buffer[58]<<0)-(layer_in_buffer[58]<<2)-(layer_in_buffer[58]<<4)-(layer_in_buffer[58]<<7)+(layer_in_buffer[58]<<11)+(layer_in_buffer[58]<<13)+(layer_in_buffer[58]<<14))-(0+(layer_in_buffer[59]<<8)+(layer_in_buffer[59]<<9)+(layer_in_buffer[59]<<12)+(layer_in_buffer[59]<<14))-(0+(layer_in_buffer[60]<<3)-(layer_in_buffer[60]<<5)-(layer_in_buffer[60]<<8)+(layer_in_buffer[60]<<11)+(layer_in_buffer[60]<<13))+(0-(layer_in_buffer[61]<<3)+(layer_in_buffer[61]<<8)+(layer_in_buffer[61]<<10)+(layer_in_buffer[61]<<11))-(0+(layer_in_buffer[62]<<6)-(layer_in_buffer[62]<<9)+(layer_in_buffer[62]<<14))-(0+(layer_in_buffer[63]<<0)+(layer_in_buffer[63]<<4)-(layer_in_buffer[63]<<7)+(layer_in_buffer[63]<<10));
wire [DATA_WIDTH-1:0]   weight_bias0;
assign weight_bias0=in_buffer_weight0+(-830);
wire [DATA_WIDTH-1:0]   weight_bias1;
assign weight_bias1=in_buffer_weight1+(-996);
wire [DATA_WIDTH-1:0]   weight_bias2;
assign weight_bias2=in_buffer_weight2+(747);
wire [DATA_WIDTH-1:0]   weight_bias3;
assign weight_bias3=in_buffer_weight3+(3154);
wire [DATA_WIDTH-1:0]   weight_bias4;
assign weight_bias4=in_buffer_weight4+(-2490);
wire [DATA_WIDTH-1:0]   weight_bias5;
assign weight_bias5=in_buffer_weight5+(1328);
wire [DATA_WIDTH-1:0]   weight_bias6;
assign weight_bias6=in_buffer_weight6+(-664);
wire [DATA_WIDTH-1:0]   weight_bias7;
assign weight_bias7=in_buffer_weight7+(2905);
wire [DATA_WIDTH-1:0]   weight_bias8;
assign weight_bias8=in_buffer_weight8+(-332);
wire [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias9=in_buffer_weight9+(0);
assign layer_out={
            weight_bias9,
            weight_bias8,
            weight_bias7,
            weight_bias6,
            weight_bias5,
            weight_bias4,
            weight_bias3,
            weight_bias2,
            weight_bias1,
            weight_bias0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule
