module layer1_cnn_144_25x64x10
(
    input clk,
    input rst,
    input [1728-1:0] layer_in,
    input valid,
    output  reg ready,
    output [36*10-1:0] layer_out
);
parameter DATA_WIDTH = 36;
parameter INPUT_DATA_CNT   =   64;
reg    signed [27-1:0]  in_buffer[0:INPUT_DATA_CNT-1];
genvar j;
generate
for(j=0;j<INPUT_DATA_CNT;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=layer_in[j*27+26:j*27+0];
                    end
            end
    end
endgenerate
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=$signed(in_buffer[0]*(-2))+$signed(in_buffer[1]*(41))+$signed(in_buffer[2]*(-27))+$signed(in_buffer[3]*(35))+$signed(in_buffer[4]*(77))+$signed(in_buffer[5]*(68))+$signed(in_buffer[6]*(-23))+$signed(in_buffer[7]*(-6))+$signed(in_buffer[8]*(-133))+$signed(in_buffer[9]*(83))+$signed(in_buffer[10]*(-20))+$signed(in_buffer[11]*(75))+$signed(in_buffer[12]*(-47))+$signed(in_buffer[13]*(-10))+$signed(in_buffer[14]*(37))+$signed(in_buffer[15]*(-133))+$signed(in_buffer[16]*(20))+$signed(in_buffer[17]*(-22))+$signed(in_buffer[18]*(-65))+$signed(in_buffer[19]*(-5))+$signed(in_buffer[20]*(4))+$signed(in_buffer[21]*(-103))+$signed(in_buffer[22]*(25))+$signed(in_buffer[23]*(-103))+$signed(in_buffer[24]*(33))+$signed(in_buffer[25]*(-32))+$signed(in_buffer[26]*(58))+$signed(in_buffer[27]*(-221))+$signed(in_buffer[28]*(-34))+$signed(in_buffer[29]*(136))+$signed(in_buffer[30]*(0))+$signed(in_buffer[31]*(24))+$signed(in_buffer[32]*(11))+$signed(in_buffer[33]*(13))+$signed(in_buffer[34]*(34))+$signed(in_buffer[35]*(2))+$signed(in_buffer[36]*(-104))+$signed(in_buffer[37]*(0))+$signed(in_buffer[38]*(15))+$signed(in_buffer[39]*(-18))+$signed(in_buffer[40]*(-6))+$signed(in_buffer[41]*(11))+$signed(in_buffer[42]*(-60))+$signed(in_buffer[43]*(1))+$signed(in_buffer[44]*(-106))+$signed(in_buffer[45]*(38))+$signed(in_buffer[46]*(14))+$signed(in_buffer[47]*(7))+$signed(in_buffer[48]*(-3))+$signed(in_buffer[49]*(96))+$signed(in_buffer[50]*(20))+$signed(in_buffer[51]*(-1))+$signed(in_buffer[52]*(1))+$signed(in_buffer[53]*(26))+$signed(in_buffer[54]*(7))+$signed(in_buffer[55]*(-97))+$signed(in_buffer[56]*(-95))+$signed(in_buffer[57]*(-58))+$signed(in_buffer[58]*(46))+$signed(in_buffer[59]*(-59))+$signed(in_buffer[60]*(0))+$signed(in_buffer[61]*(25))+$signed(in_buffer[62]*(7))+$signed(in_buffer[63]*(2));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=$signed(in_buffer[0]*(88))+$signed(in_buffer[1]*(40))+$signed(in_buffer[2]*(32))+$signed(in_buffer[3]*(-206))+$signed(in_buffer[4]*(106))+$signed(in_buffer[5]*(-89))+$signed(in_buffer[6]*(36))+$signed(in_buffer[7]*(32))+$signed(in_buffer[8]*(13))+$signed(in_buffer[9]*(-59))+$signed(in_buffer[10]*(-31))+$signed(in_buffer[11]*(43))+$signed(in_buffer[12]*(-48))+$signed(in_buffer[13]*(-32))+$signed(in_buffer[14]*(34))+$signed(in_buffer[15]*(30))+$signed(in_buffer[16]*(-57))+$signed(in_buffer[17]*(21))+$signed(in_buffer[18]*(-180))+$signed(in_buffer[19]*(0))+$signed(in_buffer[20]*(4))+$signed(in_buffer[21]*(-26))+$signed(in_buffer[22]*(-51))+$signed(in_buffer[23]*(93))+$signed(in_buffer[24]*(38))+$signed(in_buffer[25]*(-111))+$signed(in_buffer[26]*(4))+$signed(in_buffer[27]*(43))+$signed(in_buffer[28]*(44))+$signed(in_buffer[29]*(-5))+$signed(in_buffer[30]*(61))+$signed(in_buffer[31]*(30))+$signed(in_buffer[32]*(-3))+$signed(in_buffer[33]*(47))+$signed(in_buffer[34]*(-88))+$signed(in_buffer[35]*(56))+$signed(in_buffer[36]*(-13))+$signed(in_buffer[37]*(-48))+$signed(in_buffer[38]*(-18))+$signed(in_buffer[39]*(43))+$signed(in_buffer[40]*(0))+$signed(in_buffer[41]*(72))+$signed(in_buffer[42]*(142))+$signed(in_buffer[43]*(-7))+$signed(in_buffer[44]*(28))+$signed(in_buffer[45]*(-5))+$signed(in_buffer[46]*(63))+$signed(in_buffer[47]*(-98))+$signed(in_buffer[48]*(3))+$signed(in_buffer[49]*(18))+$signed(in_buffer[50]*(-168))+$signed(in_buffer[51]*(40))+$signed(in_buffer[52]*(47))+$signed(in_buffer[53]*(6))+$signed(in_buffer[54]*(-8))+$signed(in_buffer[55]*(12))+$signed(in_buffer[56]*(-9))+$signed(in_buffer[57]*(32))+$signed(in_buffer[58]*(-93))+$signed(in_buffer[59]*(-1))+$signed(in_buffer[60]*(5))+$signed(in_buffer[61]*(16))+$signed(in_buffer[62]*(-6))+$signed(in_buffer[63]*(-30));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=$signed(in_buffer[0]*(0))+$signed(in_buffer[1]*(11))+$signed(in_buffer[2]*(-4))+$signed(in_buffer[3]*(-43))+$signed(in_buffer[4]*(-4))+$signed(in_buffer[5]*(39))+$signed(in_buffer[6]*(-19))+$signed(in_buffer[7]*(56))+$signed(in_buffer[8]*(95))+$signed(in_buffer[9]*(-135))+$signed(in_buffer[10]*(21))+$signed(in_buffer[11]*(75))+$signed(in_buffer[12]*(-94))+$signed(in_buffer[13]*(-39))+$signed(in_buffer[14]*(44))+$signed(in_buffer[15]*(-190))+$signed(in_buffer[16]*(18))+$signed(in_buffer[17]*(0))+$signed(in_buffer[18]*(48))+$signed(in_buffer[19]*(-3))+$signed(in_buffer[20]*(-2))+$signed(in_buffer[21]*(-83))+$signed(in_buffer[22]*(36))+$signed(in_buffer[23]*(20))+$signed(in_buffer[24]*(51))+$signed(in_buffer[25]*(-30))+$signed(in_buffer[26]*(101))+$signed(in_buffer[27]*(-51))+$signed(in_buffer[28]*(-4))+$signed(in_buffer[29]*(-113))+$signed(in_buffer[30]*(7))+$signed(in_buffer[31]*(11))+$signed(in_buffer[32]*(13))+$signed(in_buffer[33]*(40))+$signed(in_buffer[34]*(-3))+$signed(in_buffer[35]*(74))+$signed(in_buffer[36]*(-12))+$signed(in_buffer[37]*(-36))+$signed(in_buffer[38]*(8))+$signed(in_buffer[39]*(-44))+$signed(in_buffer[40]*(15))+$signed(in_buffer[41]*(-26))+$signed(in_buffer[42]*(-6))+$signed(in_buffer[43]*(67))+$signed(in_buffer[44]*(2))+$signed(in_buffer[45]*(18))+$signed(in_buffer[46]*(28))+$signed(in_buffer[47]*(13))+$signed(in_buffer[48]*(-14))+$signed(in_buffer[49]*(103))+$signed(in_buffer[50]*(-67))+$signed(in_buffer[51]*(9))+$signed(in_buffer[52]*(-12))+$signed(in_buffer[53]*(-100))+$signed(in_buffer[54]*(-4))+$signed(in_buffer[55]*(2))+$signed(in_buffer[56]*(12))+$signed(in_buffer[57]*(60))+$signed(in_buffer[58]*(-83))+$signed(in_buffer[59]*(23))+$signed(in_buffer[60]*(-3))+$signed(in_buffer[61]*(16))+$signed(in_buffer[62]*(-16))+$signed(in_buffer[63]*(0));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=$signed(in_buffer[0]*(37))+$signed(in_buffer[1]*(33))+$signed(in_buffer[2]*(28))+$signed(in_buffer[3]*(2))+$signed(in_buffer[4]*(13))+$signed(in_buffer[5]*(-18))+$signed(in_buffer[6]*(33))+$signed(in_buffer[7]*(49))+$signed(in_buffer[8]*(-10))+$signed(in_buffer[9]*(-34))+$signed(in_buffer[10]*(2))+$signed(in_buffer[11]*(6))+$signed(in_buffer[12]*(-40))+$signed(in_buffer[13]*(0))+$signed(in_buffer[14]*(-68))+$signed(in_buffer[15]*(-9))+$signed(in_buffer[16]*(11))+$signed(in_buffer[17]*(16))+$signed(in_buffer[18]*(9))+$signed(in_buffer[19]*(0))+$signed(in_buffer[20]*(14))+$signed(in_buffer[21]*(80))+$signed(in_buffer[22]*(21))+$signed(in_buffer[23]*(6))+$signed(in_buffer[24]*(-55))+$signed(in_buffer[25]*(-2))+$signed(in_buffer[26]*(10))+$signed(in_buffer[27]*(-74))+$signed(in_buffer[28]*(61))+$signed(in_buffer[29]*(-68))+$signed(in_buffer[30]*(-59))+$signed(in_buffer[31]*(15))+$signed(in_buffer[32]*(-3))+$signed(in_buffer[33]*(-53))+$signed(in_buffer[34]*(-5))+$signed(in_buffer[35]*(-49))+$signed(in_buffer[36]*(-19))+$signed(in_buffer[37]*(24))+$signed(in_buffer[38]*(-15))+$signed(in_buffer[39]*(-79))+$signed(in_buffer[40]*(3))+$signed(in_buffer[41]*(-29))+$signed(in_buffer[42]*(89))+$signed(in_buffer[43]*(39))+$signed(in_buffer[44]*(47))+$signed(in_buffer[45]*(-27))+$signed(in_buffer[46]*(-91))+$signed(in_buffer[47]*(-18))+$signed(in_buffer[48]*(-4))+$signed(in_buffer[49]*(-27))+$signed(in_buffer[50]*(-28))+$signed(in_buffer[51]*(-16))+$signed(in_buffer[52]*(-10))+$signed(in_buffer[53]*(35))+$signed(in_buffer[54]*(8))+$signed(in_buffer[55]*(28))+$signed(in_buffer[56]*(-13))+$signed(in_buffer[57]*(-143))+$signed(in_buffer[58]*(-11))+$signed(in_buffer[59]*(16))+$signed(in_buffer[60]*(17))+$signed(in_buffer[61]*(-72))+$signed(in_buffer[62]*(-10))+$signed(in_buffer[63]*(-22));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=$signed(in_buffer[0]*(-41))+$signed(in_buffer[1]*(-147))+$signed(in_buffer[2]*(-29))+$signed(in_buffer[3]*(-2))+$signed(in_buffer[4]*(-8))+$signed(in_buffer[5]*(-101))+$signed(in_buffer[6]*(-60))+$signed(in_buffer[7]*(7))+$signed(in_buffer[8]*(15))+$signed(in_buffer[9]*(-23))+$signed(in_buffer[10]*(35))+$signed(in_buffer[11]*(-59))+$signed(in_buffer[12]*(36))+$signed(in_buffer[13]*(-46))+$signed(in_buffer[14]*(36))+$signed(in_buffer[15]*(39))+$signed(in_buffer[16]*(-16))+$signed(in_buffer[17]*(-28))+$signed(in_buffer[18]*(12))+$signed(in_buffer[19]*(-17))+$signed(in_buffer[20]*(10))+$signed(in_buffer[21]*(-13))+$signed(in_buffer[22]*(-167))+$signed(in_buffer[23]*(90))+$signed(in_buffer[24]*(-30))+$signed(in_buffer[25]*(32))+$signed(in_buffer[26]*(-84))+$signed(in_buffer[27]*(11))+$signed(in_buffer[28]*(39))+$signed(in_buffer[29]*(9))+$signed(in_buffer[30]*(-30))+$signed(in_buffer[31]*(-12))+$signed(in_buffer[32]*(-4))+$signed(in_buffer[33]*(99))+$signed(in_buffer[34]*(-13))+$signed(in_buffer[35]*(46))+$signed(in_buffer[36]*(82))+$signed(in_buffer[37]*(-47))+$signed(in_buffer[38]*(-103))+$signed(in_buffer[39]*(114))+$signed(in_buffer[40]*(0))+$signed(in_buffer[41]*(16))+$signed(in_buffer[42]*(2))+$signed(in_buffer[43]*(-13))+$signed(in_buffer[44]*(16))+$signed(in_buffer[45]*(-109))+$signed(in_buffer[46]*(-43))+$signed(in_buffer[47]*(55))+$signed(in_buffer[48]*(4))+$signed(in_buffer[49]*(-15))+$signed(in_buffer[50]*(-47))+$signed(in_buffer[51]*(-39))+$signed(in_buffer[52]*(62))+$signed(in_buffer[53]*(22))+$signed(in_buffer[54]*(4))+$signed(in_buffer[55]*(39))+$signed(in_buffer[56]*(32))+$signed(in_buffer[57]*(-43))+$signed(in_buffer[58]*(-66))+$signed(in_buffer[59]*(-65))+$signed(in_buffer[60]*(-29))+$signed(in_buffer[61]*(8))+$signed(in_buffer[62]*(-10))+$signed(in_buffer[63]*(42));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=$signed(in_buffer[0]*(33))+$signed(in_buffer[1]*(61))+$signed(in_buffer[2]*(2))+$signed(in_buffer[3]*(20))+$signed(in_buffer[4]*(-39))+$signed(in_buffer[5]*(-63))+$signed(in_buffer[6]*(98))+$signed(in_buffer[7]*(7))+$signed(in_buffer[8]*(-2))+$signed(in_buffer[9]*(70))+$signed(in_buffer[10]*(0))+$signed(in_buffer[11]*(-47))+$signed(in_buffer[12]*(71))+$signed(in_buffer[13]*(27))+$signed(in_buffer[14]*(-71))+$signed(in_buffer[15]*(89))+$signed(in_buffer[16]*(7))+$signed(in_buffer[17]*(-6))+$signed(in_buffer[18]*(68))+$signed(in_buffer[19]*(-14))+$signed(in_buffer[20]*(4))+$signed(in_buffer[21]*(105))+$signed(in_buffer[22]*(30))+$signed(in_buffer[23]*(-15))+$signed(in_buffer[24]*(-94))+$signed(in_buffer[25]*(-18))+$signed(in_buffer[26]*(79))+$signed(in_buffer[27]*(46))+$signed(in_buffer[28]*(-49))+$signed(in_buffer[29]*(-43))+$signed(in_buffer[30]*(-39))+$signed(in_buffer[31]*(18))+$signed(in_buffer[32]*(2))+$signed(in_buffer[33]*(-72))+$signed(in_buffer[34]*(10))+$signed(in_buffer[35]*(-187))+$signed(in_buffer[36]*(-150))+$signed(in_buffer[37]*(-17))+$signed(in_buffer[38]*(-33))+$signed(in_buffer[39]*(36))+$signed(in_buffer[40]*(-15))+$signed(in_buffer[41]*(-1))+$signed(in_buffer[42]*(-165))+$signed(in_buffer[43]*(-85))+$signed(in_buffer[44]*(-66))+$signed(in_buffer[45]*(40))+$signed(in_buffer[46]*(-69))+$signed(in_buffer[47]*(-9))+$signed(in_buffer[48]*(4))+$signed(in_buffer[49]*(-78))+$signed(in_buffer[50]*(36))+$signed(in_buffer[51]*(24))+$signed(in_buffer[52]*(-9))+$signed(in_buffer[53]*(26))+$signed(in_buffer[54]*(-10))+$signed(in_buffer[55]*(51))+$signed(in_buffer[56]*(-1))+$signed(in_buffer[57]*(13))+$signed(in_buffer[58]*(-1))+$signed(in_buffer[59]*(-6))+$signed(in_buffer[60]*(-19))+$signed(in_buffer[61]*(1))+$signed(in_buffer[62]*(-19))+$signed(in_buffer[63]*(-53));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=$signed(in_buffer[0]*(-4))+$signed(in_buffer[1]*(-77))+$signed(in_buffer[2]*(-53))+$signed(in_buffer[3]*(-17))+$signed(in_buffer[4]*(18))+$signed(in_buffer[5]*(-108))+$signed(in_buffer[6]*(78))+$signed(in_buffer[7]*(-106))+$signed(in_buffer[8]*(-106))+$signed(in_buffer[9]*(55))+$signed(in_buffer[10]*(1))+$signed(in_buffer[11]*(57))+$signed(in_buffer[12]*(-46))+$signed(in_buffer[13]*(-29))+$signed(in_buffer[14]*(-17))+$signed(in_buffer[15]*(-68))+$signed(in_buffer[16]*(8))+$signed(in_buffer[17]*(7))+$signed(in_buffer[18]*(67))+$signed(in_buffer[19]*(9))+$signed(in_buffer[20]*(-9))+$signed(in_buffer[21]*(-6))+$signed(in_buffer[22]*(-134))+$signed(in_buffer[23]*(-35))+$signed(in_buffer[24]*(5))+$signed(in_buffer[25]*(28))+$signed(in_buffer[26]*(35))+$signed(in_buffer[27]*(90))+$signed(in_buffer[28]*(-103))+$signed(in_buffer[29]*(74))+$signed(in_buffer[30]*(148))+$signed(in_buffer[31]*(7))+$signed(in_buffer[32]*(-1))+$signed(in_buffer[33]*(-88))+$signed(in_buffer[34]*(29))+$signed(in_buffer[35]*(-62))+$signed(in_buffer[36]*(-129))+$signed(in_buffer[37]*(25))+$signed(in_buffer[38]*(17))+$signed(in_buffer[39]*(40))+$signed(in_buffer[40]*(-10))+$signed(in_buffer[41]*(-20))+$signed(in_buffer[42]*(-94))+$signed(in_buffer[43]*(-38))+$signed(in_buffer[44]*(-70))+$signed(in_buffer[45]*(29))+$signed(in_buffer[46]*(75))+$signed(in_buffer[47]*(29))+$signed(in_buffer[48]*(-12))+$signed(in_buffer[49]*(53))+$signed(in_buffer[50]*(8))+$signed(in_buffer[51]*(-62))+$signed(in_buffer[52]*(71))+$signed(in_buffer[53]*(-27))+$signed(in_buffer[54]*(0))+$signed(in_buffer[55]*(-138))+$signed(in_buffer[56]*(-27))+$signed(in_buffer[57]*(39))+$signed(in_buffer[58]*(68))+$signed(in_buffer[59]*(19))+$signed(in_buffer[60]*(37))+$signed(in_buffer[61]*(-9))+$signed(in_buffer[62]*(12))+$signed(in_buffer[63]*(-13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=$signed(in_buffer[0]*(-14))+$signed(in_buffer[1]*(-59))+$signed(in_buffer[2]*(75))+$signed(in_buffer[3]*(-17))+$signed(in_buffer[4]*(45))+$signed(in_buffer[5]*(108))+$signed(in_buffer[6]*(-167))+$signed(in_buffer[7]*(-23))+$signed(in_buffer[8]*(9))+$signed(in_buffer[9]*(-24))+$signed(in_buffer[10]*(-26))+$signed(in_buffer[11]*(-25))+$signed(in_buffer[12]*(27))+$signed(in_buffer[13]*(24))+$signed(in_buffer[14]*(95))+$signed(in_buffer[15]*(22))+$signed(in_buffer[16]*(-63))+$signed(in_buffer[17]*(-74))+$signed(in_buffer[18]*(-100))+$signed(in_buffer[19]*(-14))+$signed(in_buffer[20]*(10))+$signed(in_buffer[21]*(-160))+$signed(in_buffer[22]*(55))+$signed(in_buffer[23]*(-12))+$signed(in_buffer[24]*(8))+$signed(in_buffer[25]*(-13))+$signed(in_buffer[26]*(-66))+$signed(in_buffer[27]*(31))+$signed(in_buffer[28]*(-5))+$signed(in_buffer[29]*(4))+$signed(in_buffer[30]*(16))+$signed(in_buffer[31]*(4))+$signed(in_buffer[32]*(11))+$signed(in_buffer[33]*(52))+$signed(in_buffer[34]*(-59))+$signed(in_buffer[35]*(-19))+$signed(in_buffer[36]*(61))+$signed(in_buffer[37]*(-18))+$signed(in_buffer[38]*(4))+$signed(in_buffer[39]*(-68))+$signed(in_buffer[40]*(14))+$signed(in_buffer[41]*(36))+$signed(in_buffer[42]*(57))+$signed(in_buffer[43]*(-61))+$signed(in_buffer[44]*(35))+$signed(in_buffer[45]*(-112))+$signed(in_buffer[46]*(-73))+$signed(in_buffer[47]*(31))+$signed(in_buffer[48]*(6))+$signed(in_buffer[49]*(-41))+$signed(in_buffer[50]*(11))+$signed(in_buffer[51]*(121))+$signed(in_buffer[52]*(-55))+$signed(in_buffer[53]*(-1))+$signed(in_buffer[54]*(-3))+$signed(in_buffer[55]*(25))+$signed(in_buffer[56]*(14))+$signed(in_buffer[57]*(-100))+$signed(in_buffer[58]*(162))+$signed(in_buffer[59]*(160))+$signed(in_buffer[60]*(-37))+$signed(in_buffer[61]*(-26))+$signed(in_buffer[62]*(-1))+$signed(in_buffer[63]*(24));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=$signed(in_buffer[0]*(-134))+$signed(in_buffer[1]*(15))+$signed(in_buffer[2]*(-3))+$signed(in_buffer[3]*(2))+$signed(in_buffer[4]*(-68))+$signed(in_buffer[5]*(-15))+$signed(in_buffer[6]*(-53))+$signed(in_buffer[7]*(4))+$signed(in_buffer[8]*(60))+$signed(in_buffer[9]*(0))+$signed(in_buffer[10]*(7))+$signed(in_buffer[11]*(-74))+$signed(in_buffer[12]*(27))+$signed(in_buffer[13]*(34))+$signed(in_buffer[14]*(-96))+$signed(in_buffer[15]*(15))+$signed(in_buffer[16]*(12))+$signed(in_buffer[17]*(6))+$signed(in_buffer[18]*(-89))+$signed(in_buffer[19]*(7))+$signed(in_buffer[20]*(-13))+$signed(in_buffer[21]*(26))+$signed(in_buffer[22]*(2))+$signed(in_buffer[23]*(-63))+$signed(in_buffer[24]*(29))+$signed(in_buffer[25]*(36))+$signed(in_buffer[26]*(-11))+$signed(in_buffer[27]*(-2))+$signed(in_buffer[28]*(-29))+$signed(in_buffer[29]*(-20))+$signed(in_buffer[30]*(48))+$signed(in_buffer[31]*(-4))+$signed(in_buffer[32]*(9))+$signed(in_buffer[33]*(-38))+$signed(in_buffer[34]*(-7))+$signed(in_buffer[35]*(-20))+$signed(in_buffer[36]*(-129))+$signed(in_buffer[37]*(20))+$signed(in_buffer[38]*(13))+$signed(in_buffer[39]*(3))+$signed(in_buffer[40]*(11))+$signed(in_buffer[41]*(-55))+$signed(in_buffer[42]*(-81))+$signed(in_buffer[43]*(-15))+$signed(in_buffer[44]*(29))+$signed(in_buffer[45]*(18))+$signed(in_buffer[46]*(30))+$signed(in_buffer[47]*(-21))+$signed(in_buffer[48]*(-18))+$signed(in_buffer[49]*(15))+$signed(in_buffer[50]*(39))+$signed(in_buffer[51]*(-91))+$signed(in_buffer[52]*(-66))+$signed(in_buffer[53]*(1))+$signed(in_buffer[54]*(-18))+$signed(in_buffer[55]*(-35))+$signed(in_buffer[56]*(16))+$signed(in_buffer[57]*(17))+$signed(in_buffer[58]*(-112))+$signed(in_buffer[59]*(3))+$signed(in_buffer[60]*(40))+$signed(in_buffer[61]*(1))+$signed(in_buffer[62]*(-6))+$signed(in_buffer[63]*(6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=$signed(in_buffer[0]*(84))+$signed(in_buffer[1]*(-31))+$signed(in_buffer[2]*(-6))+$signed(in_buffer[3]*(22))+$signed(in_buffer[4]*(-60))+$signed(in_buffer[5]*(6))+$signed(in_buffer[6]*(-123))+$signed(in_buffer[7]*(-31))+$signed(in_buffer[8]*(5))+$signed(in_buffer[9]*(14))+$signed(in_buffer[10]*(35))+$signed(in_buffer[11]*(57))+$signed(in_buffer[12]*(-6))+$signed(in_buffer[13]*(32))+$signed(in_buffer[14]*(14))+$signed(in_buffer[15]*(16))+$signed(in_buffer[16]*(5))+$signed(in_buffer[17]*(-41))+$signed(in_buffer[18]*(-22))+$signed(in_buffer[19]*(5))+$signed(in_buffer[20]*(-3))+$signed(in_buffer[21]*(3))+$signed(in_buffer[22]*(10))+$signed(in_buffer[23]*(-166))+$signed(in_buffer[24]*(-100))+$signed(in_buffer[25]*(29))+$signed(in_buffer[26]*(-134))+$signed(in_buffer[27]*(-26))+$signed(in_buffer[28]*(25))+$signed(in_buffer[29]*(27))+$signed(in_buffer[30]*(-102))+$signed(in_buffer[31]*(-62))+$signed(in_buffer[32]*(10))+$signed(in_buffer[33]*(-49))+$signed(in_buffer[34]*(-22))+$signed(in_buffer[35]*(72))+$signed(in_buffer[36]*(73))+$signed(in_buffer[37]*(23))+$signed(in_buffer[38]*(13))+$signed(in_buffer[39]*(-82))+$signed(in_buffer[40]*(14))+$signed(in_buffer[41]*(-8))+$signed(in_buffer[42]*(-2))+$signed(in_buffer[43]*(40))+$signed(in_buffer[44]*(13))+$signed(in_buffer[45]*(-10))+$signed(in_buffer[46]*(32))+$signed(in_buffer[47]*(4))+$signed(in_buffer[48]*(-14))+$signed(in_buffer[49]*(-133))+$signed(in_buffer[50]*(38))+$signed(in_buffer[51]*(-99))+$signed(in_buffer[52]*(-88))+$signed(in_buffer[53]*(20))+$signed(in_buffer[54]*(-16))+$signed(in_buffer[55]*(4))+$signed(in_buffer[56]*(40))+$signed(in_buffer[57]*(86))+$signed(in_buffer[58]*(-15))+$signed(in_buffer[59]*(-215))+$signed(in_buffer[60]*(13))+$signed(in_buffer[61]*(68))+$signed(in_buffer[62]*(9))+$signed(in_buffer[63]*(9));
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias0=in_buffer_weight0+(-82);
assign weight_bias1=in_buffer_weight1+(-23);
assign weight_bias2=in_buffer_weight2+(27);
assign weight_bias3=in_buffer_weight3+(30);
assign weight_bias4=in_buffer_weight4+(-2);
assign weight_bias5=in_buffer_weight5+(66);
assign weight_bias6=in_buffer_weight6+(-35);
assign weight_bias7=in_buffer_weight7+(21);
assign weight_bias8=in_buffer_weight8+(-21);
assign weight_bias9=in_buffer_weight9+(-6);
assign layer_out={weight_bias9,weight_bias8,weight_bias7,weight_bias6,weight_bias5,weight_bias4,weight_bias3,weight_bias2,weight_bias1,weight_bias0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule