module layer0_tcb_121x32x10
(
    input clk,
    input rst,
    input [121*8-1:0] img,
    input valid,
    output  reg ready,
    output [25*32-1:0] layer_out
);
parameter DATA_WIDTH = 25;
parameter IMG_SZ   =   121;
reg    signed [8-1:0]  in_buffer[0:IMG_SZ-1];
integer i;
always@(posedge clk )
    begin
        if(rst)
            begin
                for(i=0;i<IMG_SZ;i=i+1)
                    begin
                        in_buffer[i]<=0;
                    end
            end
        else
        begin
       in_buffer[0]<=img[7:0];
       in_buffer[1]<=img[15:8];
       in_buffer[2]<=img[23:16];
       in_buffer[3]<=img[31:24];
       in_buffer[4]<=img[39:32];
       in_buffer[5]<=img[47:40];
       in_buffer[6]<=img[55:48];
       in_buffer[7]<=img[63:56];
       in_buffer[8]<=img[71:64];
       in_buffer[9]<=img[79:72];
       in_buffer[10]<=img[87:80];
       in_buffer[11]<=img[95:88];
       in_buffer[12]<=img[103:96];
       in_buffer[13]<=img[111:104];
       in_buffer[14]<=img[119:112];
       in_buffer[15]<=img[127:120];
       in_buffer[16]<=img[135:128];
       in_buffer[17]<=img[143:136];
       in_buffer[18]<=img[151:144];
       in_buffer[19]<=img[159:152];
       in_buffer[20]<=img[167:160];
       in_buffer[21]<=img[175:168];
       in_buffer[22]<=img[183:176];
       in_buffer[23]<=img[191:184];
       in_buffer[24]<=img[199:192];
       in_buffer[25]<=img[207:200];
       in_buffer[26]<=img[215:208];
       in_buffer[27]<=img[223:216];
       in_buffer[28]<=img[231:224];
       in_buffer[29]<=img[239:232];
       in_buffer[30]<=img[247:240];
       in_buffer[31]<=img[255:248];
       in_buffer[32]<=img[263:256];
       in_buffer[33]<=img[271:264];
       in_buffer[34]<=img[279:272];
       in_buffer[35]<=img[287:280];
       in_buffer[36]<=img[295:288];
       in_buffer[37]<=img[303:296];
       in_buffer[38]<=img[311:304];
       in_buffer[39]<=img[319:312];
       in_buffer[40]<=img[327:320];
       in_buffer[41]<=img[335:328];
       in_buffer[42]<=img[343:336];
       in_buffer[43]<=img[351:344];
       in_buffer[44]<=img[359:352];
       in_buffer[45]<=img[367:360];
       in_buffer[46]<=img[375:368];
       in_buffer[47]<=img[383:376];
       in_buffer[48]<=img[391:384];
       in_buffer[49]<=img[399:392];
       in_buffer[50]<=img[407:400];
       in_buffer[51]<=img[415:408];
       in_buffer[52]<=img[423:416];
       in_buffer[53]<=img[431:424];
       in_buffer[54]<=img[439:432];
       in_buffer[55]<=img[447:440];
       in_buffer[56]<=img[455:448];
       in_buffer[57]<=img[463:456];
       in_buffer[58]<=img[471:464];
       in_buffer[59]<=img[479:472];
       in_buffer[60]<=img[487:480];
       in_buffer[61]<=img[495:488];
       in_buffer[62]<=img[503:496];
       in_buffer[63]<=img[511:504];
       in_buffer[64]<=img[519:512];
       in_buffer[65]<=img[527:520];
       in_buffer[66]<=img[535:528];
       in_buffer[67]<=img[543:536];
       in_buffer[68]<=img[551:544];
       in_buffer[69]<=img[559:552];
       in_buffer[70]<=img[567:560];
       in_buffer[71]<=img[575:568];
       in_buffer[72]<=img[583:576];
       in_buffer[73]<=img[591:584];
       in_buffer[74]<=img[599:592];
       in_buffer[75]<=img[607:600];
       in_buffer[76]<=img[615:608];
       in_buffer[77]<=img[623:616];
       in_buffer[78]<=img[631:624];
       in_buffer[79]<=img[639:632];
       in_buffer[80]<=img[647:640];
       in_buffer[81]<=img[655:648];
       in_buffer[82]<=img[663:656];
       in_buffer[83]<=img[671:664];
       in_buffer[84]<=img[679:672];
       in_buffer[85]<=img[687:680];
       in_buffer[86]<=img[695:688];
       in_buffer[87]<=img[703:696];
       in_buffer[88]<=img[711:704];
       in_buffer[89]<=img[719:712];
       in_buffer[90]<=img[727:720];
       in_buffer[91]<=img[735:728];
       in_buffer[92]<=img[743:736];
       in_buffer[93]<=img[751:744];
       in_buffer[94]<=img[759:752];
       in_buffer[95]<=img[767:760];
       in_buffer[96]<=img[775:768];
       in_buffer[97]<=img[783:776];
       in_buffer[98]<=img[791:784];
       in_buffer[99]<=img[799:792];
       in_buffer[100]<=img[807:800];
       in_buffer[101]<=img[815:808];
       in_buffer[102]<=img[823:816];
       in_buffer[103]<=img[831:824];
       in_buffer[104]<=img[839:832];
       in_buffer[105]<=img[847:840];
       in_buffer[106]<=img[855:848];
       in_buffer[107]<=img[863:856];
       in_buffer[108]<=img[871:864];
       in_buffer[109]<=img[879:872];
       in_buffer[110]<=img[887:880];
       in_buffer[111]<=img[895:888];
       in_buffer[112]<=img[903:896];
       in_buffer[113]<=img[911:904];
       in_buffer[114]<=img[919:912];
       in_buffer[115]<=img[927:920];
       in_buffer[116]<=img[935:928];
       in_buffer[117]<=img[943:936];
       in_buffer[118]<=img[951:944];
       in_buffer[119]<=img[959:952];
       in_buffer[120]<=img[967:960];
        end
   end
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0+(0+(in_buffer[0]<<5)+(in_buffer[0]<<6)+(in_buffer[0]<<9)+(in_buffer[0]<<11))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<1)-(in_buffer[1]<<4)-(in_buffer[1]<<6)-(in_buffer[1]<<8)+(in_buffer[1]<<10)+(in_buffer[1]<<11))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<3)+(in_buffer[2]<<7)+(in_buffer[2]<<12))-(0+(in_buffer[3]<<0)-(in_buffer[3]<<2)-(in_buffer[3]<<4)+(in_buffer[3]<<7)+(in_buffer[3]<<10)+(in_buffer[3]<<12))-(0-(in_buffer[4]<<2)-(in_buffer[4]<<5)+(in_buffer[4]<<8)+(in_buffer[4]<<12))+(0+(in_buffer[5]<<1)-(in_buffer[5]<<4)-(in_buffer[5]<<6)-(in_buffer[5]<<8)+(in_buffer[5]<<11)+(in_buffer[5]<<12))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<1)-(in_buffer[6]<<7)+(in_buffer[6]<<9)+(in_buffer[6]<<10))-(0+(in_buffer[7]<<0)-(in_buffer[7]<<2)+(in_buffer[7]<<5)+(in_buffer[7]<<7)+(in_buffer[7]<<8)+(in_buffer[7]<<11)+(in_buffer[7]<<12))+(0-(in_buffer[8]<<1)-(in_buffer[8]<<3)-(in_buffer[8]<<5)+(in_buffer[8]<<9)+(in_buffer[8]<<10))+(0+(in_buffer[9]<<0)-(in_buffer[9]<<2)+(in_buffer[9]<<5)+(in_buffer[9]<<7)+(in_buffer[9]<<8)+(in_buffer[9]<<11)+(in_buffer[9]<<12))+(0-(in_buffer[10]<<1)-(in_buffer[10]<<4)-(in_buffer[10]<<7)-(in_buffer[10]<<10)+(in_buffer[10]<<13)+(in_buffer[10]<<14))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<4)+(in_buffer[11]<<7)+(in_buffer[11]<<9)+(in_buffer[11]<<11)+(in_buffer[11]<<14))+(0+(in_buffer[12]<<2)+(in_buffer[12]<<3)+(in_buffer[12]<<6)+(in_buffer[12]<<8))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<4)-(in_buffer[13]<<6)-(in_buffer[13]<<8)+(in_buffer[13]<<11))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<3)+(in_buffer[14]<<5)+(in_buffer[14]<<9)+(in_buffer[14]<<10))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<5)+(in_buffer[15]<<7)+(in_buffer[15]<<8))+(0-(in_buffer[16]<<4)+(in_buffer[16]<<9)+(in_buffer[16]<<11)+(in_buffer[16]<<12))-(0+(in_buffer[17]<<0)-(in_buffer[17]<<3)+(in_buffer[17]<<8))+(0-(in_buffer[18]<<0)-(in_buffer[18]<<3)+(in_buffer[18]<<6)+(in_buffer[18]<<10))-(0+(in_buffer[19]<<0)-(in_buffer[19]<<3)+(in_buffer[19]<<8))+(0-(in_buffer[20]<<3)-(in_buffer[20]<<6)+(in_buffer[20]<<9)+(in_buffer[20]<<13))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<5)+(in_buffer[21]<<7)+(in_buffer[21]<<10)+(in_buffer[21]<<12)+(in_buffer[21]<<14))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<2)+(in_buffer[22]<<4)+(in_buffer[22]<<7)+(in_buffer[22]<<9)+(in_buffer[22]<<10)+(in_buffer[22]<<13))-(0-(in_buffer[24]<<0)+(in_buffer[24]<<4)+(in_buffer[24]<<5)+(in_buffer[24]<<8)+(in_buffer[24]<<12))-(0+(in_buffer[25]<<1)+(in_buffer[25]<<3)+(in_buffer[25]<<6)+(in_buffer[25]<<8)+(in_buffer[25]<<11)+(in_buffer[25]<<12))-(0-(in_buffer[26]<<0)+(in_buffer[26]<<5)+(in_buffer[26]<<6)-(in_buffer[26]<<9)+(in_buffer[26]<<11)+(in_buffer[26]<<12))+(0+(in_buffer[27]<<1)+(in_buffer[27]<<5)-(in_buffer[27]<<8)+(in_buffer[27]<<11))-(0-(in_buffer[28]<<0)+(in_buffer[28]<<3)+(in_buffer[28]<<4)+(in_buffer[28]<<7)-(in_buffer[28]<<9)+(in_buffer[28]<<12))-(0-(in_buffer[29]<<0)+(in_buffer[29]<<4)+(in_buffer[29]<<5)+(in_buffer[29]<<8)+(in_buffer[29]<<12))-(0+(in_buffer[30]<<0)-(in_buffer[30]<<3)-(in_buffer[30]<<5)-(in_buffer[30]<<7)+(in_buffer[30]<<10)+(in_buffer[30]<<11))+(0-(in_buffer[31]<<1)-(in_buffer[31]<<3)+(in_buffer[31]<<6)+(in_buffer[31]<<12))+(0-(in_buffer[32]<<1)+(in_buffer[32]<<6)+(in_buffer[32]<<7)-(in_buffer[32]<<10)+(in_buffer[32]<<12)+(in_buffer[32]<<13))+(0+(in_buffer[33]<<1)+(in_buffer[33]<<3)+(in_buffer[33]<<6)+(in_buffer[33]<<8)+(in_buffer[33]<<11)+(in_buffer[33]<<12))+(0-(in_buffer[34]<<0)+(in_buffer[34]<<4)-(in_buffer[34]<<6)-(in_buffer[34]<<8)+(in_buffer[34]<<11))-(0-(in_buffer[35]<<0)-(in_buffer[35]<<3)+(in_buffer[35]<<6)+(in_buffer[35]<<10))+(0-(in_buffer[36]<<0)+(in_buffer[36]<<3)-(in_buffer[36]<<6)+(in_buffer[36]<<10)+(in_buffer[36]<<12))-(0-(in_buffer[37]<<0)+(in_buffer[37]<<3)-(in_buffer[37]<<5)+(in_buffer[37]<<7)+(in_buffer[37]<<8)+(in_buffer[37]<<11))-(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)-(in_buffer[38]<<4)+(in_buffer[38]<<8)+(in_buffer[38]<<9))-(0-(in_buffer[39]<<0)+(in_buffer[39]<<4)-(in_buffer[39]<<6)-(in_buffer[39]<<8)+(in_buffer[39]<<11))+(0-(in_buffer[40]<<0)+(in_buffer[40]<<2)+(in_buffer[40]<<3)+(in_buffer[40]<<6)+(in_buffer[40]<<8)+(in_buffer[40]<<10)+(in_buffer[40]<<11))+(0-(in_buffer[41]<<2)+(in_buffer[41]<<7)+(in_buffer[41]<<9)+(in_buffer[41]<<10))+(0-(in_buffer[42]<<1)-(in_buffer[42]<<3)+(in_buffer[42]<<6)+(in_buffer[42]<<12))+(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6)-(in_buffer[43]<<8)+(in_buffer[43]<<11)+(in_buffer[43]<<13))+(0+(in_buffer[44]<<1)+(in_buffer[44]<<3)+(in_buffer[44]<<7)+(in_buffer[44]<<10))-(0+(in_buffer[45]<<0)+(in_buffer[45]<<1)+(in_buffer[45]<<4)+(in_buffer[45]<<6))-(0+(in_buffer[46]<<1)-(in_buffer[46]<<3)-(in_buffer[46]<<6)+(in_buffer[46]<<9)+(in_buffer[46]<<11))+(0+(in_buffer[47]<<0)-(in_buffer[47]<<2)-(in_buffer[47]<<4)+(in_buffer[47]<<7)+(in_buffer[47]<<10)+(in_buffer[47]<<12))-(0+(in_buffer[48]<<1)+(in_buffer[48]<<3)+(in_buffer[48]<<4)+(in_buffer[48]<<10)+(in_buffer[48]<<12))-(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)-(in_buffer[49]<<4)+(in_buffer[49]<<8)+(in_buffer[49]<<9))+(0+(in_buffer[50]<<3)+(in_buffer[50]<<4)+(in_buffer[50]<<7)+(in_buffer[50]<<9))+(0+(in_buffer[51]<<1)+(in_buffer[51]<<3)+(in_buffer[51]<<5)-(in_buffer[51]<<7)+(in_buffer[51]<<10)+(in_buffer[51]<<13))-(0+(in_buffer[52]<<2)+(in_buffer[52]<<3)+(in_buffer[52]<<6)+(in_buffer[52]<<8))+(0+(in_buffer[53]<<0)+(in_buffer[53]<<2)-(in_buffer[53]<<4)-(in_buffer[53]<<7)+(in_buffer[53]<<11))+(0-(in_buffer[54]<<0)-(in_buffer[54]<<2)-(in_buffer[54]<<4)-(in_buffer[54]<<6)+(in_buffer[54]<<11)+(in_buffer[54]<<12))-(0+(in_buffer[55]<<0)+(in_buffer[55]<<5)+(in_buffer[55]<<8)+(in_buffer[55]<<9)+(in_buffer[55]<<12))-(0+(in_buffer[56]<<1)+(in_buffer[56]<<5)-(in_buffer[56]<<8)+(in_buffer[56]<<11))-(0+(in_buffer[57]<<1)+(in_buffer[57]<<3)+(in_buffer[57]<<7)+(in_buffer[57]<<10))+(0-(in_buffer[58]<<0)-(in_buffer[58]<<2)-(in_buffer[58]<<4)+(in_buffer[58]<<8)+(in_buffer[58]<<9))-(0+(in_buffer[59]<<0)-(in_buffer[59]<<3)-(in_buffer[59]<<5)-(in_buffer[59]<<7)+(in_buffer[59]<<10)+(in_buffer[59]<<11))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)-(in_buffer[60]<<4)-(in_buffer[60]<<6)-(in_buffer[60]<<8)+(in_buffer[60]<<10)+(in_buffer[60]<<11))-(0+(in_buffer[61]<<5)+(in_buffer[61]<<6)+(in_buffer[61]<<9)+(in_buffer[61]<<11))+(0+(in_buffer[62]<<0)+(in_buffer[62]<<2)+(in_buffer[62]<<5)+(in_buffer[62]<<7)+(in_buffer[62]<<10)+(in_buffer[62]<<11))-(0-(in_buffer[63]<<1)-(in_buffer[63]<<3)+(in_buffer[63]<<6)+(in_buffer[63]<<12))+(0+(in_buffer[64]<<4)+(in_buffer[64]<<5)+(in_buffer[64]<<8)+(in_buffer[64]<<10))-(0-(in_buffer[65]<<0)+(in_buffer[65]<<4)-(in_buffer[65]<<6)-(in_buffer[65]<<8)+(in_buffer[65]<<11))-(0-(in_buffer[66]<<0)+(in_buffer[66]<<4)+(in_buffer[66]<<5)+(in_buffer[66]<<8)+(in_buffer[66]<<12))+(0+(in_buffer[67]<<0)-(in_buffer[67]<<2)-(in_buffer[67]<<4)+(in_buffer[67]<<7)+(in_buffer[67]<<10)+(in_buffer[67]<<12))+(0+(in_buffer[68]<<0)+(in_buffer[68]<<2)+(in_buffer[68]<<3)+(in_buffer[68]<<9)+(in_buffer[68]<<11))-(0+(in_buffer[69]<<1)+(in_buffer[69]<<2)-(in_buffer[69]<<8)+(in_buffer[69]<<10)+(in_buffer[69]<<11))-(0+(in_buffer[70]<<0)-(in_buffer[70]<<4)-(in_buffer[70]<<9)+(in_buffer[70]<<12))-(0+(in_buffer[71]<<0)+(in_buffer[71]<<2)+(in_buffer[71]<<3)+(in_buffer[71]<<9)+(in_buffer[71]<<11))-(0-(in_buffer[72]<<0)+(in_buffer[72]<<2)+(in_buffer[72]<<3)+(in_buffer[72]<<6)+(in_buffer[72]<<8)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0+(in_buffer[73]<<0)+(in_buffer[73]<<4)-(in_buffer[73]<<7)+(in_buffer[73]<<10))-(0-(in_buffer[74]<<2)+(in_buffer[74]<<7)+(in_buffer[74]<<9)+(in_buffer[74]<<10))+(0+(in_buffer[75]<<1)+(in_buffer[75]<<4)+(in_buffer[75]<<6)+(in_buffer[75]<<10)+(in_buffer[75]<<11))+(0+(in_buffer[76]<<0)-(in_buffer[76]<<2)+(in_buffer[76]<<6)-(in_buffer[76]<<8)+(in_buffer[76]<<12))+(0-(in_buffer[77]<<2)+(in_buffer[77]<<7)+(in_buffer[77]<<9)+(in_buffer[77]<<10))+(0-(in_buffer[78]<<0)+(in_buffer[78]<<3)-(in_buffer[78]<<5)+(in_buffer[78]<<7)+(in_buffer[78]<<8)+(in_buffer[78]<<11))-(0+(in_buffer[79]<<0)+(in_buffer[79]<<2)+(in_buffer[79]<<4)-(in_buffer[79]<<6)+(in_buffer[79]<<9)+(in_buffer[79]<<12))-(0+(in_buffer[80]<<0)+(in_buffer[80]<<1)-(in_buffer[80]<<4)-(in_buffer[80]<<6)-(in_buffer[80]<<8)+(in_buffer[80]<<10)+(in_buffer[80]<<11))-(0+(in_buffer[81]<<1)-(in_buffer[81]<<4)+(in_buffer[81]<<9))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)-(in_buffer[82]<<4)+(in_buffer[82]<<8)+(in_buffer[82]<<9))+(0+(in_buffer[83]<<1)+(in_buffer[83]<<2)+(in_buffer[83]<<5)+(in_buffer[83]<<7))+(0+(in_buffer[84]<<0)-(in_buffer[84]<<3)+(in_buffer[84]<<8))-(0+(in_buffer[85]<<0)+(in_buffer[85]<<1)-(in_buffer[85]<<4)-(in_buffer[85]<<6)-(in_buffer[85]<<8)+(in_buffer[85]<<10)+(in_buffer[85]<<11))+(0+(in_buffer[86]<<0)+(in_buffer[86]<<5)+(in_buffer[86]<<8)+(in_buffer[86]<<9)+(in_buffer[86]<<12))+(0-(in_buffer[87]<<1)+(in_buffer[87]<<4)+(in_buffer[87]<<5)+(in_buffer[87]<<8)-(in_buffer[87]<<10)+(in_buffer[87]<<13))-(0+(in_buffer[88]<<0)-(in_buffer[88]<<2)-(in_buffer[88]<<5)+(in_buffer[88]<<8)+(in_buffer[88]<<10))+(0-(in_buffer[89]<<1)+(in_buffer[89]<<6)+(in_buffer[89]<<8)+(in_buffer[89]<<9))+(0-(in_buffer[90]<<2)+(in_buffer[90]<<7)+(in_buffer[90]<<9)+(in_buffer[90]<<10))+(0+(in_buffer[91]<<0)+(in_buffer[91]<<2)-(in_buffer[91]<<4)-(in_buffer[91]<<7)+(in_buffer[91]<<11))+(0-(in_buffer[92]<<0)+(in_buffer[92]<<5)+(in_buffer[92]<<7)+(in_buffer[92]<<8))+(0+(in_buffer[93]<<3)-(in_buffer[93]<<6)+(in_buffer[93]<<11))-(0-(in_buffer[94]<<0)-(in_buffer[94]<<2)+(in_buffer[94]<<5)+(in_buffer[94]<<11))-(0-(in_buffer[95]<<1)+(in_buffer[95]<<6)+(in_buffer[95]<<8)+(in_buffer[95]<<9))+(0-(in_buffer[96]<<0)+(in_buffer[96]<<4)-(in_buffer[96]<<7)-(in_buffer[96]<<10)+(in_buffer[96]<<13))+(0-(in_buffer[97]<<0)+(in_buffer[97]<<3)+(in_buffer[97]<<5)-(in_buffer[97]<<9)+(in_buffer[97]<<13))+(0-(in_buffer[98]<<1)+(in_buffer[98]<<11)+(in_buffer[98]<<12))-(0+(in_buffer[99]<<3)-(in_buffer[99]<<6)+(in_buffer[99]<<11))-(0+(in_buffer[100]<<0)+(in_buffer[100]<<4)-(in_buffer[100]<<7)+(in_buffer[100]<<10))+(0-(in_buffer[101]<<1)-(in_buffer[101]<<3)+(in_buffer[101]<<6)+(in_buffer[101]<<12))+(0+(in_buffer[102]<<1)+(in_buffer[102]<<2)-(in_buffer[102]<<5)-(in_buffer[102]<<7)-(in_buffer[102]<<9)+(in_buffer[102]<<11)+(in_buffer[102]<<12))+(0+(in_buffer[103]<<1)-(in_buffer[103]<<4)+(in_buffer[103]<<9))+(0-(in_buffer[104]<<0)+(in_buffer[104]<<4)-(in_buffer[104]<<6)-(in_buffer[104]<<8)+(in_buffer[104]<<11))-(0-(in_buffer[105]<<0)+(in_buffer[105]<<5)+(in_buffer[105]<<7)+(in_buffer[105]<<8))+(0+(in_buffer[106]<<0)+(in_buffer[106]<<3)+(in_buffer[106]<<7)+(in_buffer[106]<<12))+(0+(in_buffer[107]<<0)+(in_buffer[107]<<2)-(in_buffer[107]<<8)+(in_buffer[107]<<11)+(in_buffer[107]<<12))+(0-(in_buffer[108]<<0)-(in_buffer[108]<<3)+(in_buffer[108]<<6)+(in_buffer[108]<<10))-(0+(in_buffer[109]<<3)-(in_buffer[109]<<6)+(in_buffer[109]<<11))+(0-(in_buffer[110]<<1)-(in_buffer[110]<<3)+(in_buffer[110]<<6)+(in_buffer[110]<<12))+(0+(in_buffer[111]<<1)+(in_buffer[111]<<5)-(in_buffer[111]<<8)+(in_buffer[111]<<11))-(0+(in_buffer[112]<<2)+(in_buffer[112]<<4)+(in_buffer[112]<<8)+(in_buffer[112]<<11))+(0+(in_buffer[114]<<1)-(in_buffer[114]<<5)-(in_buffer[114]<<10)+(in_buffer[114]<<13))+(0+(in_buffer[115]<<3)-(in_buffer[115]<<5)-(in_buffer[115]<<8)+(in_buffer[115]<<11)+(in_buffer[115]<<13))+(0-(in_buffer[116]<<3)+(in_buffer[116]<<8)+(in_buffer[116]<<10)+(in_buffer[116]<<11))+(0+(in_buffer[117]<<4)-(in_buffer[117]<<7)+(in_buffer[117]<<12))-(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<5)+(in_buffer[118]<<11))-(0+(in_buffer[119]<<3)-(in_buffer[119]<<6)+(in_buffer[119]<<11))-(0+(in_buffer[120]<<0)-(in_buffer[120]<<2)+(in_buffer[120]<<10)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0-(0+(in_buffer[0]<<1)-(in_buffer[0]<<4)+(in_buffer[0]<<9))-(0-(in_buffer[1]<<2)+(in_buffer[1]<<6)+(in_buffer[1]<<7)+(in_buffer[1]<<10)+(in_buffer[1]<<14))-(0+(in_buffer[2]<<6)+(in_buffer[2]<<7)+(in_buffer[2]<<10)+(in_buffer[2]<<12))+(0+(in_buffer[3]<<2)-(in_buffer[3]<<5)-(in_buffer[3]<<7)-(in_buffer[3]<<9)+(in_buffer[3]<<12)+(in_buffer[3]<<13))+(0+(in_buffer[4]<<2)+(in_buffer[4]<<8)+(in_buffer[4]<<9)+(in_buffer[4]<<13))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3)+(in_buffer[5]<<9)+(in_buffer[5]<<13))+(0+(in_buffer[6]<<2)+(in_buffer[6]<<3)-(in_buffer[6]<<9)+(in_buffer[6]<<11)+(in_buffer[6]<<12))+(0-(in_buffer[7]<<3)+(in_buffer[7]<<7)-(in_buffer[7]<<9)-(in_buffer[7]<<11)+(in_buffer[7]<<14))+(0-(in_buffer[8]<<0)+(in_buffer[8]<<5)+(in_buffer[8]<<6)-(in_buffer[8]<<9)+(in_buffer[8]<<11)+(in_buffer[8]<<12))-(0-(in_buffer[9]<<1)-(in_buffer[9]<<3)+(in_buffer[9]<<6)+(in_buffer[9]<<12))-(0-(in_buffer[10]<<1)+(in_buffer[10]<<5)-(in_buffer[10]<<7)-(in_buffer[10]<<9)+(in_buffer[10]<<12))+(0+(in_buffer[11]<<0)-(in_buffer[11]<<3)-(in_buffer[11]<<5)-(in_buffer[11]<<7)+(in_buffer[11]<<10)+(in_buffer[11]<<11))-(0-(in_buffer[12]<<3)+(in_buffer[12]<<8)+(in_buffer[12]<<10)+(in_buffer[12]<<11))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<3)+(in_buffer[13]<<4)+(in_buffer[13]<<7)-(in_buffer[13]<<9)+(in_buffer[13]<<12))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)-(in_buffer[14]<<4)-(in_buffer[14]<<7)+(in_buffer[14]<<11))-(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<5)+(in_buffer[15]<<11))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<4)-(in_buffer[16]<<6)-(in_buffer[16]<<8)+(in_buffer[16]<<11))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<4)-(in_buffer[17]<<7)+(in_buffer[17]<<10))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)-(in_buffer[18]<<4)-(in_buffer[18]<<7)+(in_buffer[18]<<11))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<2)+(in_buffer[19]<<5)+(in_buffer[19]<<7))+(0-(in_buffer[20]<<0)-(in_buffer[20]<<2)+(in_buffer[20]<<5)+(in_buffer[20]<<7)+(in_buffer[20]<<8)+(in_buffer[20]<<12)+(in_buffer[20]<<13))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<3)-(in_buffer[21]<<5)-(in_buffer[21]<<8)+(in_buffer[21]<<12))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<2)+(in_buffer[22]<<5)+(in_buffer[22]<<9)+(in_buffer[22]<<11)+(in_buffer[22]<<13))+(0-(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<3)+(in_buffer[23]<<6)+(in_buffer[23]<<8)+(in_buffer[23]<<10)+(in_buffer[23]<<11))+(0+(in_buffer[24]<<3)-(in_buffer[24]<<6)+(in_buffer[24]<<11))-(0-(in_buffer[25]<<2)+(in_buffer[25]<<7)+(in_buffer[25]<<9)+(in_buffer[25]<<10))+(0-(in_buffer[26]<<0)-(in_buffer[26]<<3)+(in_buffer[26]<<6)+(in_buffer[26]<<10))+(0+(in_buffer[27]<<0)+(in_buffer[27]<<1)-(in_buffer[27]<<4)-(in_buffer[27]<<6)-(in_buffer[27]<<8)+(in_buffer[27]<<10)+(in_buffer[27]<<11))+(0+(in_buffer[28]<<0)+(in_buffer[28]<<1)-(in_buffer[28]<<7)+(in_buffer[28]<<9)+(in_buffer[28]<<10))+(0+(in_buffer[29]<<1)-(in_buffer[29]<<4)+(in_buffer[29]<<9))+(0+(in_buffer[30]<<0)+(in_buffer[30]<<1)+(in_buffer[30]<<4)+(in_buffer[30]<<6))+(0-(in_buffer[31]<<0)-(in_buffer[31]<<2)-(in_buffer[31]<<4)+(in_buffer[31]<<7)-(in_buffer[31]<<10)+(in_buffer[31]<<12)+(in_buffer[31]<<13))+(0-(in_buffer[32]<<3)-(in_buffer[32]<<6)+(in_buffer[32]<<9)+(in_buffer[32]<<13))+(0-(in_buffer[33]<<1)-(in_buffer[33]<<3)+(in_buffer[33]<<6)+(in_buffer[33]<<12))+(0+(in_buffer[34]<<1)+(in_buffer[34]<<3)+(in_buffer[34]<<4)+(in_buffer[34]<<10)+(in_buffer[34]<<12))+(0+(in_buffer[35]<<0)+(in_buffer[35]<<2)+(in_buffer[35]<<3)+(in_buffer[35]<<9)+(in_buffer[35]<<11))-(0+(in_buffer[36]<<0)+(in_buffer[36]<<1)-(in_buffer[36]<<7)+(in_buffer[36]<<9)+(in_buffer[36]<<10))-(0-(in_buffer[37]<<0)+(in_buffer[37]<<5)+(in_buffer[37]<<7)+(in_buffer[37]<<8))-(0+(in_buffer[38]<<1)-(in_buffer[38]<<4)+(in_buffer[38]<<9))-(0-(in_buffer[39]<<0)+(in_buffer[39]<<3)-(in_buffer[39]<<5)+(in_buffer[39]<<7)+(in_buffer[39]<<8)+(in_buffer[39]<<11))-(0+(in_buffer[40]<<1)-(in_buffer[40]<<4)+(in_buffer[40]<<9))+(0+(in_buffer[41]<<2)-(in_buffer[41]<<5)+(in_buffer[41]<<10))+(0+(in_buffer[42]<<1)+(in_buffer[42]<<3)+(in_buffer[42]<<5)-(in_buffer[42]<<7)+(in_buffer[42]<<10)+(in_buffer[42]<<13))-(0-(in_buffer[43]<<2)+(in_buffer[43]<<7)+(in_buffer[43]<<9)+(in_buffer[43]<<10))+(0+(in_buffer[44]<<0)+(in_buffer[44]<<1)-(in_buffer[44]<<4)-(in_buffer[44]<<6)-(in_buffer[44]<<8)+(in_buffer[44]<<10)+(in_buffer[44]<<11))+(0-(in_buffer[45]<<0)-(in_buffer[45]<<2)+(in_buffer[45]<<5)+(in_buffer[45]<<11))-(0+(in_buffer[46]<<0)-(in_buffer[46]<<3)+(in_buffer[46]<<8))-(0+(in_buffer[47]<<0)+(in_buffer[47]<<5)+(in_buffer[47]<<8)+(in_buffer[47]<<9)+(in_buffer[47]<<12))+(0-(in_buffer[48]<<0)-(in_buffer[48]<<2)-(in_buffer[48]<<4)+(in_buffer[48]<<8)+(in_buffer[48]<<9))-(0+(in_buffer[49]<<0)-(in_buffer[49]<<3)+(in_buffer[49]<<8))+(0-(in_buffer[50]<<0)-(in_buffer[50]<<2)+(in_buffer[50]<<5)+(in_buffer[50]<<11))-(0+(in_buffer[51]<<1)+(in_buffer[51]<<3)+(in_buffer[51]<<4)+(in_buffer[51]<<10)+(in_buffer[51]<<12))-(0-(in_buffer[52]<<2)-(in_buffer[52]<<4)-(in_buffer[52]<<6)+(in_buffer[52]<<10)+(in_buffer[52]<<11))+(0+(in_buffer[53]<<1)-(in_buffer[53]<<3)-(in_buffer[53]<<6)+(in_buffer[53]<<9)+(in_buffer[53]<<11))-(0+(in_buffer[54]<<0)+(in_buffer[54]<<2)-(in_buffer[54]<<5)+(in_buffer[54]<<7)+(in_buffer[54]<<8)+(in_buffer[54]<<13))+(0-(in_buffer[55]<<0)+(in_buffer[55]<<4)+(in_buffer[55]<<6)+(in_buffer[55]<<12)+(in_buffer[55]<<13))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<3)+(in_buffer[56]<<9)+(in_buffer[56]<<11))-(0-(in_buffer[57]<<1)-(in_buffer[57]<<3)-(in_buffer[57]<<5)+(in_buffer[57]<<9)+(in_buffer[57]<<10))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)+(in_buffer[58]<<3)+(in_buffer[58]<<9)+(in_buffer[58]<<11))+(0+(in_buffer[59]<<5)+(in_buffer[59]<<6)+(in_buffer[59]<<9)+(in_buffer[59]<<11))+(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)+(in_buffer[60]<<4)+(in_buffer[60]<<6))+(0-(in_buffer[61]<<0)+(in_buffer[61]<<10)+(in_buffer[61]<<11))-(0-(in_buffer[62]<<0)+(in_buffer[62]<<2)+(in_buffer[62]<<3)+(in_buffer[62]<<6)+(in_buffer[62]<<8)+(in_buffer[62]<<10)+(in_buffer[62]<<11))-(0-(in_buffer[63]<<0)+(in_buffer[63]<<3)+(in_buffer[63]<<5)-(in_buffer[63]<<9)+(in_buffer[63]<<13))-(0-(in_buffer[64]<<1)+(in_buffer[64]<<5)-(in_buffer[64]<<7)-(in_buffer[64]<<9)+(in_buffer[64]<<12))+(0+(in_buffer[65]<<2)-(in_buffer[65]<<5)+(in_buffer[65]<<10))-(0+(in_buffer[66]<<0)+(in_buffer[66]<<3)+(in_buffer[66]<<7)+(in_buffer[66]<<12))-(0-(in_buffer[67]<<1)+(in_buffer[67]<<6)+(in_buffer[67]<<8)+(in_buffer[67]<<9))+(0+(in_buffer[68]<<0)+(in_buffer[68]<<4)-(in_buffer[68]<<7)+(in_buffer[68]<<10))+(0+(in_buffer[69]<<0)+(in_buffer[69]<<2)-(in_buffer[69]<<4)-(in_buffer[69]<<7)+(in_buffer[69]<<11))+(0+(in_buffer[70]<<2)-(in_buffer[70]<<4)-(in_buffer[70]<<7)+(in_buffer[70]<<10)+(in_buffer[70]<<12))-(0+(in_buffer[71]<<0)+(in_buffer[71]<<1)+(in_buffer[71]<<4)+(in_buffer[71]<<6))+(0-(in_buffer[72]<<0)+(in_buffer[72]<<4)+(in_buffer[72]<<5)+(in_buffer[72]<<8)+(in_buffer[72]<<12))-(0-(in_buffer[73]<<1)-(in_buffer[73]<<3)-(in_buffer[73]<<5)+(in_buffer[73]<<9)+(in_buffer[73]<<10))-(0+(in_buffer[74]<<0)+(in_buffer[74]<<1)+(in_buffer[74]<<6)+(in_buffer[74]<<9)+(in_buffer[74]<<11)+(in_buffer[74]<<12))-(0+(in_buffer[75]<<0)+(in_buffer[75]<<2)+(in_buffer[75]<<3)+(in_buffer[75]<<9)+(in_buffer[75]<<11))-(0-(in_buffer[77]<<1)-(in_buffer[77]<<4)-(in_buffer[77]<<7)-(in_buffer[77]<<10)+(in_buffer[77]<<13)+(in_buffer[77]<<14))-(0+(in_buffer[78]<<1)+(in_buffer[78]<<3)+(in_buffer[78]<<4)+(in_buffer[78]<<10)+(in_buffer[78]<<12))+(0+(in_buffer[79]<<2)+(in_buffer[79]<<3)+(in_buffer[79]<<6)+(in_buffer[79]<<8))+(0-(in_buffer[80]<<0)+(in_buffer[80]<<4)+(in_buffer[80]<<5)+(in_buffer[80]<<8)+(in_buffer[80]<<12))+(0+(in_buffer[81]<<1)-(in_buffer[81]<<4)-(in_buffer[81]<<6)-(in_buffer[81]<<8)+(in_buffer[81]<<11)+(in_buffer[81]<<12))-(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)-(in_buffer[82]<<4)+(in_buffer[82]<<8)+(in_buffer[82]<<9))+(0+(in_buffer[83]<<2)+(in_buffer[83]<<6)-(in_buffer[83]<<9)+(in_buffer[83]<<12))+(0+(in_buffer[84]<<0)+(in_buffer[84]<<1)+(in_buffer[84]<<4)+(in_buffer[84]<<8)+(in_buffer[84]<<10)+(in_buffer[84]<<12))-(0-(in_buffer[85]<<1)+(in_buffer[85]<<11)+(in_buffer[85]<<12))-(0-(in_buffer[86]<<1)-(in_buffer[86]<<3)+(in_buffer[86]<<8)+(in_buffer[86]<<10)+(in_buffer[86]<<13))-(0-(in_buffer[87]<<0)+(in_buffer[87]<<2)+(in_buffer[87]<<3)+(in_buffer[87]<<9)+(in_buffer[87]<<13))-(0-(in_buffer[88]<<1)-(in_buffer[88]<<3)-(in_buffer[88]<<5)+(in_buffer[88]<<8)-(in_buffer[88]<<11)+(in_buffer[88]<<13)+(in_buffer[88]<<14))-(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)-(in_buffer[89]<<10)+(in_buffer[89]<<14))-(0-(in_buffer[90]<<1)+(in_buffer[90]<<11)+(in_buffer[90]<<12))+(0-(in_buffer[91]<<1)-(in_buffer[91]<<3)+(in_buffer[91]<<6)+(in_buffer[91]<<12))+(0+(in_buffer[92]<<0)+(in_buffer[92]<<2)-(in_buffer[92]<<8)+(in_buffer[92]<<11)+(in_buffer[92]<<12))-(0+(in_buffer[93]<<0)+(in_buffer[93]<<2)-(in_buffer[93]<<4)-(in_buffer[93]<<7)+(in_buffer[93]<<11))+(0+(in_buffer[94]<<5)+(in_buffer[94]<<6)+(in_buffer[94]<<9)+(in_buffer[94]<<11))+(0+(in_buffer[95]<<1)+(in_buffer[95]<<3)-(in_buffer[95]<<5)-(in_buffer[95]<<8)+(in_buffer[95]<<12))-(0+(in_buffer[96]<<2)+(in_buffer[96]<<4)-(in_buffer[96]<<6)-(in_buffer[96]<<9)+(in_buffer[96]<<13))-(0+(in_buffer[97]<<0)+(in_buffer[97]<<2)+(in_buffer[97]<<6)+(in_buffer[97]<<8)+(in_buffer[97]<<10)+(in_buffer[97]<<12)+(in_buffer[97]<<14))-(0-(in_buffer[98]<<0)-(in_buffer[98]<<2)+(in_buffer[98]<<6)-(in_buffer[98]<<8)+(in_buffer[98]<<11)+(in_buffer[98]<<13))-(0-(in_buffer[99]<<2)-(in_buffer[99]<<5)+(in_buffer[99]<<10)+(in_buffer[99]<<13)+(in_buffer[99]<<14))-(0-(in_buffer[100]<<0)+(in_buffer[100]<<4)-(in_buffer[100]<<7)-(in_buffer[100]<<10)+(in_buffer[100]<<13))+(0+(in_buffer[101]<<4)+(in_buffer[101]<<5)+(in_buffer[101]<<8)+(in_buffer[101]<<10))+(0+(in_buffer[102]<<1)+(in_buffer[102]<<4)+(in_buffer[102]<<6)+(in_buffer[102]<<10)+(in_buffer[102]<<11))-(0-(in_buffer[103]<<0)-(in_buffer[103]<<2)-(in_buffer[103]<<4)+(in_buffer[103]<<8)+(in_buffer[103]<<9))-(0+(in_buffer[104]<<2)+(in_buffer[104]<<3)-(in_buffer[104]<<9)+(in_buffer[104]<<11)+(in_buffer[104]<<12))+(0+(in_buffer[105]<<2)+(in_buffer[105]<<3)+(in_buffer[105]<<6)+(in_buffer[105]<<8))+(0+(in_buffer[106]<<2)+(in_buffer[106]<<4)+(in_buffer[106]<<8)+(in_buffer[106]<<11))-(0+(in_buffer[107]<<0)+(in_buffer[107]<<1)-(in_buffer[107]<<4)-(in_buffer[107]<<6)-(in_buffer[107]<<8)+(in_buffer[107]<<10)+(in_buffer[107]<<11))-(0+(in_buffer[108]<<0)+(in_buffer[108]<<4)-(in_buffer[108]<<6)+(in_buffer[108]<<9)+(in_buffer[108]<<14))-(0+(in_buffer[109]<<0)-(in_buffer[109]<<3)+(in_buffer[109]<<6)+(in_buffer[109]<<7)+(in_buffer[109]<<11)+(in_buffer[109]<<13)+(in_buffer[109]<<14))-(0+(in_buffer[110]<<1)-(in_buffer[110]<<3)+(in_buffer[110]<<5)+(in_buffer[110]<<6)+(in_buffer[110]<<9)+(in_buffer[110]<<12)+(in_buffer[110]<<14))+(0+(in_buffer[111]<<0)+(in_buffer[111]<<3)+(in_buffer[111]<<5)+(in_buffer[111]<<9)+(in_buffer[111]<<10))+(0-(in_buffer[112]<<2)+(in_buffer[112]<<7)+(in_buffer[112]<<9)+(in_buffer[112]<<10))+(0-(in_buffer[113]<<3)-(in_buffer[113]<<5)-(in_buffer[113]<<7)+(in_buffer[113]<<11)+(in_buffer[113]<<12))-(0-(in_buffer[114]<<1)+(in_buffer[114]<<6)+(in_buffer[114]<<8)+(in_buffer[114]<<9))-(0+(in_buffer[115]<<0)-(in_buffer[115]<<2)-(in_buffer[115]<<4)+(in_buffer[115]<<7)+(in_buffer[115]<<10)+(in_buffer[115]<<12))-(0+(in_buffer[116]<<4)+(in_buffer[116]<<5)+(in_buffer[116]<<8)+(in_buffer[116]<<10))+(0-(in_buffer[117]<<1)-(in_buffer[117]<<3)+(in_buffer[117]<<6)+(in_buffer[117]<<12))-(0+(in_buffer[119]<<1)+(in_buffer[119]<<2)+(in_buffer[119]<<5)+(in_buffer[119]<<7))-(0-(in_buffer[120]<<0)+(in_buffer[120]<<3)+(in_buffer[120]<<7)+(in_buffer[120]<<11)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0-(0+(in_buffer[0]<<2)+(in_buffer[0]<<3)+(in_buffer[0]<<6)+(in_buffer[0]<<8))-(0+(in_buffer[1]<<2)+(in_buffer[1]<<3)+(in_buffer[1]<<6)+(in_buffer[1]<<8))+(0+(in_buffer[2]<<6)+(in_buffer[2]<<7)+(in_buffer[2]<<10)+(in_buffer[2]<<12))+(0+(in_buffer[3]<<1)-(in_buffer[3]<<4)+(in_buffer[3]<<9))-(0-(in_buffer[4]<<0)-(in_buffer[4]<<3)-(in_buffer[4]<<5)-(in_buffer[4]<<7)+(in_buffer[4]<<10)+(in_buffer[4]<<13))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<7)+(in_buffer[5]<<11)+(in_buffer[5]<<13))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<3)-(in_buffer[6]<<5)-(in_buffer[6]<<8)-(in_buffer[6]<<10)+(in_buffer[6]<<13))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<7)+(in_buffer[7]<<12))+(0-(in_buffer[8]<<1)-(in_buffer[8]<<4)+(in_buffer[8]<<7)+(in_buffer[8]<<11))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<3)+(in_buffer[9]<<6)+(in_buffer[9]<<8)+(in_buffer[9]<<11)+(in_buffer[9]<<12))+(0+(in_buffer[10]<<2)+(in_buffer[10]<<3)+(in_buffer[10]<<6)+(in_buffer[10]<<10)+(in_buffer[10]<<12)+(in_buffer[10]<<14))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<3)-(in_buffer[11]<<5)+(in_buffer[11]<<7)+(in_buffer[11]<<8)+(in_buffer[11]<<11))-(0+(in_buffer[12]<<3)+(in_buffer[12]<<5)+(in_buffer[12]<<9)+(in_buffer[12]<<12))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<3)+(in_buffer[13]<<7)+(in_buffer[13]<<12))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<6)+(in_buffer[14]<<7)+(in_buffer[14]<<11))-(0-(in_buffer[15]<<1)+(in_buffer[15]<<6)+(in_buffer[15]<<8)+(in_buffer[15]<<9))-(0+(in_buffer[16]<<3)+(in_buffer[16]<<4)+(in_buffer[16]<<7)+(in_buffer[16]<<9))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<3)+(in_buffer[17]<<9)+(in_buffer[17]<<11))-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)-(in_buffer[18]<<4)+(in_buffer[18]<<8)+(in_buffer[18]<<9))-(0+(in_buffer[19]<<1)-(in_buffer[19]<<4)-(in_buffer[19]<<6)-(in_buffer[19]<<8)+(in_buffer[19]<<11)+(in_buffer[19]<<12))-(0-(in_buffer[20]<<0)+(in_buffer[20]<<5)+(in_buffer[20]<<7)+(in_buffer[20]<<8))+(0-(in_buffer[21]<<5)+(in_buffer[21]<<10)+(in_buffer[21]<<12)+(in_buffer[21]<<13))+(0-(in_buffer[22]<<0)+(in_buffer[22]<<3)+(in_buffer[22]<<7)+(in_buffer[22]<<11)+(in_buffer[22]<<13))-(0+(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<4)+(in_buffer[23]<<5)+(in_buffer[23]<<8)+(in_buffer[23]<<11)+(in_buffer[23]<<13))-(0-(in_buffer[24]<<2)+(in_buffer[24]<<6)-(in_buffer[24]<<8)-(in_buffer[24]<<10)+(in_buffer[24]<<13))+(0-(in_buffer[25]<<1)+(in_buffer[25]<<6)+(in_buffer[25]<<8)+(in_buffer[25]<<9))-(0-(in_buffer[26]<<4)+(in_buffer[26]<<9)+(in_buffer[26]<<11)+(in_buffer[26]<<12))-(0+(in_buffer[27]<<1)+(in_buffer[27]<<7)+(in_buffer[27]<<8)+(in_buffer[27]<<12))-(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)+(in_buffer[28]<<7)+(in_buffer[28]<<9)+(in_buffer[28]<<12))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<1)-(in_buffer[29]<<7)+(in_buffer[29]<<9)+(in_buffer[29]<<10))-(0+(in_buffer[30]<<0)+(in_buffer[30]<<1)+(in_buffer[30]<<4)+(in_buffer[30]<<8)+(in_buffer[30]<<10)+(in_buffer[30]<<12))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<4)+(in_buffer[31]<<6)+(in_buffer[31]<<11)+(in_buffer[31]<<12))+(0+(in_buffer[32]<<0)+(in_buffer[32]<<4)+(in_buffer[32]<<8)-(in_buffer[32]<<10)+(in_buffer[32]<<12)+(in_buffer[32]<<13))+(0+(in_buffer[33]<<1)+(in_buffer[33]<<4)+(in_buffer[33]<<8)+(in_buffer[33]<<13))-(0+(in_buffer[34]<<2)+(in_buffer[34]<<5)+(in_buffer[34]<<7)+(in_buffer[34]<<11)+(in_buffer[34]<<12))-(0+(in_buffer[35]<<0)+(in_buffer[35]<<5)+(in_buffer[35]<<8)+(in_buffer[35]<<9)+(in_buffer[35]<<12))+(0+(in_buffer[36]<<0)+(in_buffer[36]<<5)+(in_buffer[36]<<8)+(in_buffer[36]<<9)+(in_buffer[36]<<12))-(0-(in_buffer[37]<<2)-(in_buffer[37]<<4)-(in_buffer[37]<<6)+(in_buffer[37]<<10)+(in_buffer[37]<<11))-(0-(in_buffer[38]<<2)+(in_buffer[38]<<7)+(in_buffer[38]<<9)+(in_buffer[38]<<10))+(0-(in_buffer[39]<<1)-(in_buffer[39]<<4)+(in_buffer[39]<<7)+(in_buffer[39]<<11))+(0+(in_buffer[40]<<1)-(in_buffer[40]<<4)-(in_buffer[40]<<6)-(in_buffer[40]<<8)+(in_buffer[40]<<11)+(in_buffer[40]<<12))-(0+(in_buffer[41]<<5)+(in_buffer[41]<<6)+(in_buffer[41]<<9)+(in_buffer[41]<<11))-(0-(in_buffer[42]<<1)-(in_buffer[42]<<4)+(in_buffer[42]<<7)+(in_buffer[42]<<11))+(0-(in_buffer[43]<<1)+(in_buffer[43]<<11)+(in_buffer[43]<<12))+(0-(in_buffer[44]<<2)-(in_buffer[44]<<4)-(in_buffer[44]<<6)+(in_buffer[44]<<10)+(in_buffer[44]<<11))-(0-(in_buffer[45]<<0)+(in_buffer[45]<<4)-(in_buffer[45]<<6)-(in_buffer[45]<<8)+(in_buffer[45]<<11))-(0+(in_buffer[46]<<0)+(in_buffer[46]<<1)-(in_buffer[46]<<4)-(in_buffer[46]<<6)-(in_buffer[46]<<8)+(in_buffer[46]<<10)+(in_buffer[46]<<11))+(0+(in_buffer[47]<<1)+(in_buffer[47]<<3)+(in_buffer[47]<<7)+(in_buffer[47]<<10))-(0+(in_buffer[48]<<0)+(in_buffer[48]<<1)+(in_buffer[48]<<4)+(in_buffer[48]<<6))+(0+(in_buffer[49]<<1)-(in_buffer[49]<<4)+(in_buffer[49]<<9))+(0+(in_buffer[50]<<3)-(in_buffer[50]<<6)+(in_buffer[50]<<11))+(0+(in_buffer[51]<<0)+(in_buffer[51]<<1)+(in_buffer[51]<<4)+(in_buffer[51]<<8)+(in_buffer[51]<<10)+(in_buffer[51]<<12))+(0+(in_buffer[52]<<0)-(in_buffer[52]<<2)-(in_buffer[52]<<5)+(in_buffer[52]<<8)+(in_buffer[52]<<10))+(0-(in_buffer[53]<<0)+(in_buffer[53]<<3)-(in_buffer[53]<<5)+(in_buffer[53]<<7)+(in_buffer[53]<<8)+(in_buffer[53]<<11))-(0-(in_buffer[54]<<1)-(in_buffer[54]<<3)-(in_buffer[54]<<5)+(in_buffer[54]<<9)+(in_buffer[54]<<10))+(0+(in_buffer[55]<<2)+(in_buffer[55]<<3)+(in_buffer[55]<<6)+(in_buffer[55]<<8))-(0+(in_buffer[56]<<1)+(in_buffer[56]<<3)+(in_buffer[56]<<7)+(in_buffer[56]<<10))-(0-(in_buffer[57]<<1)-(in_buffer[57]<<3)-(in_buffer[57]<<5)+(in_buffer[57]<<9)+(in_buffer[57]<<10))-(0+(in_buffer[58]<<0)-(in_buffer[58]<<2)-(in_buffer[58]<<5)+(in_buffer[58]<<8)+(in_buffer[58]<<10))+(0+(in_buffer[59]<<2)+(in_buffer[59]<<4)+(in_buffer[59]<<8)+(in_buffer[59]<<11))+(0-(in_buffer[60]<<0)+(in_buffer[60]<<3)-(in_buffer[60]<<5)+(in_buffer[60]<<7)+(in_buffer[60]<<8)+(in_buffer[60]<<11))+(0-(in_buffer[61]<<0)+(in_buffer[61]<<10)+(in_buffer[61]<<11))+(0+(in_buffer[62]<<1)+(in_buffer[62]<<3)-(in_buffer[62]<<5)-(in_buffer[62]<<8)+(in_buffer[62]<<12))+(0+(in_buffer[63]<<1)+(in_buffer[63]<<3)+(in_buffer[63]<<7)+(in_buffer[63]<<10))-(0+(in_buffer[64]<<2)+(in_buffer[64]<<3)+(in_buffer[64]<<6)+(in_buffer[64]<<8))-(0+(in_buffer[65]<<1)-(in_buffer[65]<<5)-(in_buffer[65]<<10)+(in_buffer[65]<<13))+(0+(in_buffer[66]<<2)-(in_buffer[66]<<5)+(in_buffer[66]<<10))+(0+(in_buffer[67]<<0)-(in_buffer[67]<<3)-(in_buffer[67]<<6)-(in_buffer[67]<<9)+(in_buffer[67]<<11)+(in_buffer[67]<<12))+(0+(in_buffer[68]<<1)-(in_buffer[68]<<3)-(in_buffer[68]<<6)+(in_buffer[68]<<9)+(in_buffer[68]<<11))-(0+(in_buffer[69]<<2)-(in_buffer[69]<<5)+(in_buffer[69]<<10))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<2)-(in_buffer[70]<<4)-(in_buffer[70]<<7)+(in_buffer[70]<<11))+(0+(in_buffer[71]<<2)+(in_buffer[71]<<6)-(in_buffer[71]<<9)+(in_buffer[71]<<12))+(0+(in_buffer[72]<<0)+(in_buffer[72]<<2)+(in_buffer[72]<<5)+(in_buffer[72]<<7)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0+(in_buffer[73]<<0)+(in_buffer[73]<<1)-(in_buffer[73]<<7)+(in_buffer[73]<<9)+(in_buffer[73]<<10))+(0+(in_buffer[74]<<0)+(in_buffer[74]<<2)-(in_buffer[74]<<4)-(in_buffer[74]<<7)+(in_buffer[74]<<11))+(0+(in_buffer[75]<<0)+(in_buffer[75]<<1)-(in_buffer[75]<<4)-(in_buffer[75]<<6)-(in_buffer[75]<<8)+(in_buffer[75]<<10)+(in_buffer[75]<<11))-(0+(in_buffer[76]<<1)-(in_buffer[76]<<3)+(in_buffer[76]<<7)-(in_buffer[76]<<9)+(in_buffer[76]<<13))-(0+(in_buffer[77]<<3)+(in_buffer[77]<<5)+(in_buffer[77]<<9)+(in_buffer[77]<<12))+(0+(in_buffer[78]<<1)-(in_buffer[78]<<4)-(in_buffer[78]<<6)-(in_buffer[78]<<8)+(in_buffer[78]<<11)+(in_buffer[78]<<12))+(0+(in_buffer[79]<<0)+(in_buffer[79]<<1)+(in_buffer[79]<<4)+(in_buffer[79]<<6))+(0-(in_buffer[80]<<1)-(in_buffer[80]<<3)-(in_buffer[80]<<5)+(in_buffer[80]<<9)+(in_buffer[80]<<10))+(0-(in_buffer[81]<<2)+(in_buffer[81]<<7)+(in_buffer[81]<<9)+(in_buffer[81]<<10))+(0+(in_buffer[82]<<0)+(in_buffer[82]<<2)-(in_buffer[82]<<4)-(in_buffer[82]<<7)+(in_buffer[82]<<11))-(0+(in_buffer[83]<<1)-(in_buffer[83]<<4)+(in_buffer[83]<<9))+(0+(in_buffer[84]<<1)+(in_buffer[84]<<4)+(in_buffer[84]<<6)+(in_buffer[84]<<10)+(in_buffer[84]<<11))+(0-(in_buffer[85]<<1)+(in_buffer[85]<<5)-(in_buffer[85]<<7)-(in_buffer[85]<<9)+(in_buffer[85]<<12))+(0+(in_buffer[86]<<0)+(in_buffer[86]<<2)+(in_buffer[86]<<4)-(in_buffer[86]<<6)+(in_buffer[86]<<9)+(in_buffer[86]<<12))-(0+(in_buffer[87]<<0)+(in_buffer[87]<<6)+(in_buffer[87]<<7)+(in_buffer[87]<<11))-(0+(in_buffer[88]<<0)+(in_buffer[88]<<2)+(in_buffer[88]<<3)+(in_buffer[88]<<9)+(in_buffer[88]<<11))+(0+(in_buffer[89]<<0)+(in_buffer[89]<<3)+(in_buffer[89]<<4)+(in_buffer[89]<<13))+(0+(in_buffer[90]<<2)+(in_buffer[90]<<6)-(in_buffer[90]<<9)+(in_buffer[90]<<12))+(0+(in_buffer[91]<<2)+(in_buffer[91]<<5)+(in_buffer[91]<<7)+(in_buffer[91]<<11)+(in_buffer[91]<<12))+(0+(in_buffer[92]<<0)+(in_buffer[92]<<2)+(in_buffer[92]<<3)+(in_buffer[92]<<9)+(in_buffer[92]<<11))+(0+(in_buffer[93]<<0)+(in_buffer[93]<<1)-(in_buffer[93]<<7)+(in_buffer[93]<<9)+(in_buffer[93]<<10))-(0+(in_buffer[94]<<0)+(in_buffer[94]<<4)-(in_buffer[94]<<7)+(in_buffer[94]<<10))+(0+(in_buffer[95]<<0)-(in_buffer[95]<<2)+(in_buffer[95]<<6)-(in_buffer[95]<<8)+(in_buffer[95]<<12))+(0+(in_buffer[96]<<2)+(in_buffer[96]<<4)-(in_buffer[96]<<6)-(in_buffer[96]<<9)+(in_buffer[96]<<13))+(0+(in_buffer[97]<<1)+(in_buffer[97]<<3)-(in_buffer[97]<<5)-(in_buffer[97]<<8)+(in_buffer[97]<<12))+(0-(in_buffer[99]<<1)+(in_buffer[99]<<5)-(in_buffer[99]<<7)-(in_buffer[99]<<9)+(in_buffer[99]<<12))+(0+(in_buffer[100]<<2)+(in_buffer[100]<<4)+(in_buffer[100]<<8)+(in_buffer[100]<<11))+(0-(in_buffer[101]<<2)-(in_buffer[101]<<5)+(in_buffer[101]<<8)+(in_buffer[101]<<12))+(0-(in_buffer[102]<<0)+(in_buffer[102]<<4)+(in_buffer[102]<<5)+(in_buffer[102]<<8)+(in_buffer[102]<<12))+(0-(in_buffer[103]<<1)-(in_buffer[103]<<4)+(in_buffer[103]<<7)+(in_buffer[103]<<11))+(0+(in_buffer[104]<<2)+(in_buffer[104]<<4)+(in_buffer[104]<<8)+(in_buffer[104]<<11))-(0+(in_buffer[105]<<0)+(in_buffer[105]<<1)-(in_buffer[105]<<4)-(in_buffer[105]<<6)-(in_buffer[105]<<8)+(in_buffer[105]<<10)+(in_buffer[105]<<11))-(0-(in_buffer[106]<<0)+(in_buffer[106]<<3)-(in_buffer[106]<<5)+(in_buffer[106]<<7)+(in_buffer[106]<<8)+(in_buffer[106]<<11))+(0-(in_buffer[107]<<2)-(in_buffer[107]<<4)-(in_buffer[107]<<6)+(in_buffer[107]<<10)+(in_buffer[107]<<11))-(0+(in_buffer[109]<<0)+(in_buffer[109]<<2)+(in_buffer[109]<<3)+(in_buffer[109]<<9)+(in_buffer[109]<<11))-(0-(in_buffer[110]<<0)+(in_buffer[110]<<4)+(in_buffer[110]<<5)+(in_buffer[110]<<8)+(in_buffer[110]<<12))+(0+(in_buffer[111]<<3)+(in_buffer[111]<<5)+(in_buffer[111]<<9)+(in_buffer[111]<<12))+(0+(in_buffer[112]<<2)+(in_buffer[112]<<4)-(in_buffer[112]<<6)-(in_buffer[112]<<9)+(in_buffer[112]<<13))+(0+(in_buffer[113]<<5)+(in_buffer[113]<<6)+(in_buffer[113]<<9)+(in_buffer[113]<<11))+(0+(in_buffer[114]<<0)-(in_buffer[114]<<2)-(in_buffer[114]<<4)+(in_buffer[114]<<7)+(in_buffer[114]<<10)+(in_buffer[114]<<12))+(0+(in_buffer[115]<<6)+(in_buffer[115]<<7)+(in_buffer[115]<<10)+(in_buffer[115]<<12))-(0-(in_buffer[116]<<0)+(in_buffer[116]<<5)+(in_buffer[116]<<7)+(in_buffer[116]<<8))-(0-(in_buffer[117]<<2)+(in_buffer[117]<<6)-(in_buffer[117]<<8)-(in_buffer[117]<<10)+(in_buffer[117]<<13))+(0+(in_buffer[118]<<1)+(in_buffer[118]<<5)-(in_buffer[118]<<8)+(in_buffer[118]<<11))-(0+(in_buffer[119]<<0)-(in_buffer[119]<<3)+(in_buffer[119]<<8))-(0+(in_buffer[120]<<0)-(in_buffer[120]<<3)+(in_buffer[120]<<7)+(in_buffer[120]<<9)+(in_buffer[120]<<11)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0+(0+(in_buffer[0]<<1)-(in_buffer[0]<<3)-(in_buffer[0]<<6)+(in_buffer[0]<<9)+(in_buffer[0]<<11))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)-(in_buffer[1]<<5)+(in_buffer[1]<<7)+(in_buffer[1]<<8)+(in_buffer[1]<<13))-(0+(in_buffer[2]<<1)-(in_buffer[2]<<3)+(in_buffer[2]<<6)+(in_buffer[2]<<8)+(in_buffer[2]<<9)+(in_buffer[2]<<12)+(in_buffer[2]<<13))-(0-(in_buffer[3]<<1)+(in_buffer[3]<<3)+(in_buffer[3]<<4)+(in_buffer[3]<<10)+(in_buffer[3]<<14))-(0-(in_buffer[4]<<1)+(in_buffer[4]<<5)-(in_buffer[4]<<7)-(in_buffer[4]<<9)+(in_buffer[4]<<12))+(0+(in_buffer[5]<<0)-(in_buffer[5]<<4)-(in_buffer[5]<<6)+(in_buffer[5]<<8)+(in_buffer[5]<<9)+(in_buffer[5]<<13))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<4)-(in_buffer[6]<<7)+(in_buffer[6]<<10))-(0+(in_buffer[7]<<3)+(in_buffer[7]<<9)+(in_buffer[7]<<10)+(in_buffer[7]<<14))-(0+(in_buffer[8]<<1)+(in_buffer[8]<<3)+(in_buffer[8]<<5)+(in_buffer[8]<<6)-(in_buffer[8]<<11)+(in_buffer[8]<<14))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<6)+(in_buffer[9]<<9))-(0+(in_buffer[10]<<2)-(in_buffer[10]<<5)+(in_buffer[10]<<10))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<3)-(in_buffer[11]<<5)-(in_buffer[11]<<7)+(in_buffer[11]<<10)+(in_buffer[11]<<13))+(0-(in_buffer[12]<<3)-(in_buffer[12]<<5)-(in_buffer[12]<<7)+(in_buffer[12]<<11)+(in_buffer[12]<<12))+(0+(in_buffer[13]<<0)+(in_buffer[13]<<1)-(in_buffer[13]<<5)+(in_buffer[13]<<12))-(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)-(in_buffer[14]<<5)+(in_buffer[14]<<8)+(in_buffer[14]<<10))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<5)+(in_buffer[15]<<7)+(in_buffer[15]<<8))-(0-(in_buffer[16]<<1)+(in_buffer[16]<<6)+(in_buffer[16]<<8)+(in_buffer[16]<<9))+(0-(in_buffer[17]<<1)-(in_buffer[17]<<4)+(in_buffer[17]<<7)+(in_buffer[17]<<11))-(0-(in_buffer[18]<<1)-(in_buffer[18]<<3)-(in_buffer[18]<<5)+(in_buffer[18]<<9)+(in_buffer[18]<<10))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<3)-(in_buffer[19]<<5)-(in_buffer[19]<<8)+(in_buffer[19]<<12))+(0+(in_buffer[20]<<2)+(in_buffer[20]<<5)+(in_buffer[20]<<9)+(in_buffer[20]<<14))+(0-(in_buffer[21]<<0)-(in_buffer[21]<<2)-(in_buffer[21]<<4)-(in_buffer[21]<<6)+(in_buffer[21]<<11)+(in_buffer[21]<<12))+(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)-(in_buffer[22]<<4)-(in_buffer[22]<<6)+(in_buffer[22]<<11)+(in_buffer[22]<<12))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)-(in_buffer[23]<<5)+(in_buffer[23]<<12))+(0+(in_buffer[24]<<3)+(in_buffer[24]<<7)-(in_buffer[24]<<10)+(in_buffer[24]<<13))+(0-(in_buffer[25]<<0)-(in_buffer[25]<<3)+(in_buffer[25]<<6)+(in_buffer[25]<<10))-(0+(in_buffer[26]<<0)-(in_buffer[26]<<3)-(in_buffer[26]<<5)-(in_buffer[26]<<7)+(in_buffer[26]<<10)+(in_buffer[26]<<11))-(0+(in_buffer[27]<<2)+(in_buffer[27]<<5)+(in_buffer[27]<<7)+(in_buffer[27]<<11)+(in_buffer[27]<<12))-(0+(in_buffer[28]<<0)-(in_buffer[28]<<2)-(in_buffer[28]<<5)+(in_buffer[28]<<8)+(in_buffer[28]<<10))+(0-(in_buffer[29]<<1)+(in_buffer[29]<<5)-(in_buffer[29]<<7)-(in_buffer[29]<<9)+(in_buffer[29]<<12))+(0+(in_buffer[30]<<1)-(in_buffer[30]<<3)-(in_buffer[30]<<6)+(in_buffer[30]<<9)+(in_buffer[30]<<11))+(0+(in_buffer[31]<<2)+(in_buffer[31]<<5)+(in_buffer[31]<<7)+(in_buffer[31]<<11)+(in_buffer[31]<<12))+(0+(in_buffer[32]<<0)+(in_buffer[32]<<2)-(in_buffer[32]<<8)+(in_buffer[32]<<11)+(in_buffer[32]<<12))+(0-(in_buffer[33]<<3)+(in_buffer[33]<<8)+(in_buffer[33]<<10)+(in_buffer[33]<<11))+(0+(in_buffer[34]<<5)+(in_buffer[34]<<6)+(in_buffer[34]<<9)+(in_buffer[34]<<11))+(0+(in_buffer[35]<<2)+(in_buffer[35]<<4)+(in_buffer[35]<<5)+(in_buffer[35]<<11)+(in_buffer[35]<<13))+(0+(in_buffer[36]<<0)+(in_buffer[36]<<2)-(in_buffer[36]<<8)+(in_buffer[36]<<11)+(in_buffer[36]<<12))-(0+(in_buffer[37]<<0)+(in_buffer[37]<<1)-(in_buffer[37]<<5)+(in_buffer[37]<<12))-(0-(in_buffer[38]<<1)+(in_buffer[38]<<11)+(in_buffer[38]<<12))-(0-(in_buffer[39]<<0)-(in_buffer[39]<<3)+(in_buffer[39]<<6)+(in_buffer[39]<<10))+(0-(in_buffer[40]<<2)+(in_buffer[40]<<7)+(in_buffer[40]<<9)+(in_buffer[40]<<10))+(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)-(in_buffer[41]<<4)-(in_buffer[41]<<6)+(in_buffer[41]<<11)+(in_buffer[41]<<12))+(0+(in_buffer[42]<<0)+(in_buffer[42]<<2)+(in_buffer[42]<<3)+(in_buffer[42]<<9)+(in_buffer[42]<<11))+(0+(in_buffer[43]<<1)+(in_buffer[43]<<3)-(in_buffer[43]<<5)-(in_buffer[43]<<8)+(in_buffer[43]<<12))+(0+(in_buffer[44]<<1)+(in_buffer[44]<<4)+(in_buffer[44]<<6)+(in_buffer[44]<<10)+(in_buffer[44]<<11))+(0+(in_buffer[45]<<0)+(in_buffer[45]<<4)-(in_buffer[45]<<7)+(in_buffer[45]<<10))+(0-(in_buffer[46]<<0)+(in_buffer[46]<<2)+(in_buffer[46]<<3)+(in_buffer[46]<<6)+(in_buffer[46]<<8)+(in_buffer[46]<<10)+(in_buffer[46]<<11))+(0+(in_buffer[47]<<1)+(in_buffer[47]<<7)+(in_buffer[47]<<8)+(in_buffer[47]<<12))+(0+(in_buffer[48]<<0)+(in_buffer[48]<<2)+(in_buffer[48]<<6)+(in_buffer[48]<<9))-(0+(in_buffer[49]<<0)+(in_buffer[49]<<1)-(in_buffer[49]<<5)+(in_buffer[49]<<12))-(0+(in_buffer[50]<<0)-(in_buffer[50]<<3)+(in_buffer[50]<<8))+(0+(in_buffer[51]<<2)-(in_buffer[51]<<5)+(in_buffer[51]<<10))+(0+(in_buffer[52]<<1)+(in_buffer[52]<<4)+(in_buffer[52]<<6)+(in_buffer[52]<<10)+(in_buffer[52]<<11))+(0+(in_buffer[53]<<0)+(in_buffer[53]<<2)+(in_buffer[53]<<6)+(in_buffer[53]<<9))+(0+(in_buffer[54]<<1)-(in_buffer[54]<<3)-(in_buffer[54]<<6)+(in_buffer[54]<<9)+(in_buffer[54]<<11))+(0+(in_buffer[55]<<0)+(in_buffer[55]<<6)+(in_buffer[55]<<7)+(in_buffer[55]<<11))-(0-(in_buffer[56]<<2)-(in_buffer[56]<<4)-(in_buffer[56]<<6)+(in_buffer[56]<<10)+(in_buffer[56]<<11))+(0+(in_buffer[57]<<0)+(in_buffer[57]<<1)+(in_buffer[57]<<4)+(in_buffer[57]<<6))+(0-(in_buffer[58]<<1)+(in_buffer[58]<<6)+(in_buffer[58]<<8)+(in_buffer[58]<<9))-(0+(in_buffer[59]<<0)+(in_buffer[59]<<2)-(in_buffer[59]<<4)-(in_buffer[59]<<7)+(in_buffer[59]<<11))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<2)+(in_buffer[60]<<5)+(in_buffer[60]<<7)+(in_buffer[60]<<10)+(in_buffer[60]<<11))-(0-(in_buffer[61]<<0)+(in_buffer[61]<<4)-(in_buffer[61]<<6)-(in_buffer[61]<<8)+(in_buffer[61]<<11))-(0-(in_buffer[62]<<1)+(in_buffer[62]<<6)+(in_buffer[62]<<8)+(in_buffer[62]<<9))+(0+(in_buffer[64]<<0)+(in_buffer[64]<<3)+(in_buffer[64]<<5)+(in_buffer[64]<<9)+(in_buffer[64]<<10))-(0+(in_buffer[65]<<4)+(in_buffer[65]<<5)+(in_buffer[65]<<8)+(in_buffer[65]<<10))-(0+(in_buffer[66]<<0)+(in_buffer[66]<<2)+(in_buffer[66]<<4)-(in_buffer[66]<<6)+(in_buffer[66]<<9)+(in_buffer[66]<<12))-(0+(in_buffer[67]<<0)-(in_buffer[67]<<2)+(in_buffer[67]<<6)-(in_buffer[67]<<8)+(in_buffer[67]<<12))+(0+(in_buffer[68]<<0)+(in_buffer[68]<<2)+(in_buffer[68]<<3)+(in_buffer[68]<<9)+(in_buffer[68]<<11))-(0-(in_buffer[69]<<1)-(in_buffer[69]<<3)-(in_buffer[69]<<5)+(in_buffer[69]<<9)+(in_buffer[69]<<10))+(0+(in_buffer[70]<<2)-(in_buffer[70]<<5)+(in_buffer[70]<<10))+(0+(in_buffer[71]<<0)+(in_buffer[71]<<1)-(in_buffer[71]<<7)+(in_buffer[71]<<9)+(in_buffer[71]<<10))+(0+(in_buffer[72]<<2)-(in_buffer[72]<<5)+(in_buffer[72]<<10))-(0-(in_buffer[73]<<0)+(in_buffer[73]<<10)+(in_buffer[73]<<11))+(0+(in_buffer[74]<<0)+(in_buffer[74]<<1)-(in_buffer[74]<<7)+(in_buffer[74]<<9)+(in_buffer[74]<<10))+(0-(in_buffer[75]<<0)+(in_buffer[75]<<2)+(in_buffer[75]<<3)+(in_buffer[75]<<6)+(in_buffer[75]<<8)+(in_buffer[75]<<10)+(in_buffer[75]<<11))-(0-(in_buffer[76]<<1)-(in_buffer[76]<<3)+(in_buffer[76]<<6)+(in_buffer[76]<<12))+(0-(in_buffer[77]<<0)+(in_buffer[77]<<3)-(in_buffer[77]<<5)+(in_buffer[77]<<7)+(in_buffer[77]<<8)+(in_buffer[77]<<11))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<3)+(in_buffer[78]<<6)+(in_buffer[78]<<10))-(0-(in_buffer[79]<<0)-(in_buffer[79]<<2)-(in_buffer[79]<<4)+(in_buffer[79]<<8)+(in_buffer[79]<<9))-(0-(in_buffer[80]<<0)+(in_buffer[80]<<10)+(in_buffer[80]<<11))-(0+(in_buffer[81]<<1)+(in_buffer[81]<<3)+(in_buffer[81]<<7)+(in_buffer[81]<<10))+(0+(in_buffer[82]<<0)+(in_buffer[82]<<1)+(in_buffer[82]<<4)+(in_buffer[82]<<6))-(0-(in_buffer[83]<<0)+(in_buffer[83]<<5)+(in_buffer[83]<<7)+(in_buffer[83]<<8))-(0+(in_buffer[84]<<5)+(in_buffer[84]<<6)+(in_buffer[84]<<9)+(in_buffer[84]<<11))-(0-(in_buffer[85]<<1)+(in_buffer[85]<<6)+(in_buffer[85]<<8)+(in_buffer[85]<<9))+(0+(in_buffer[86]<<2)+(in_buffer[86]<<3)+(in_buffer[86]<<6)+(in_buffer[86]<<8))+(0+(in_buffer[87]<<3)-(in_buffer[87]<<6)+(in_buffer[87]<<11))+(0-(in_buffer[88]<<1)-(in_buffer[88]<<3)-(in_buffer[88]<<5)+(in_buffer[88]<<9)+(in_buffer[88]<<10))+(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<5)+(in_buffer[89]<<11))-(0+(in_buffer[90]<<0)+(in_buffer[90]<<6)+(in_buffer[90]<<7)+(in_buffer[90]<<11))-(0+(in_buffer[91]<<1)-(in_buffer[91]<<3)-(in_buffer[91]<<6)+(in_buffer[91]<<9)+(in_buffer[91]<<11))-(0-(in_buffer[92]<<0)+(in_buffer[92]<<10)+(in_buffer[92]<<11))+(0-(in_buffer[93]<<0)+(in_buffer[93]<<5)+(in_buffer[93]<<7)+(in_buffer[93]<<8))+(0+(in_buffer[94]<<0)-(in_buffer[94]<<4)-(in_buffer[94]<<9)+(in_buffer[94]<<12))+(0+(in_buffer[95]<<1)+(in_buffer[95]<<2)-(in_buffer[95]<<8)+(in_buffer[95]<<10)+(in_buffer[95]<<11))-(0-(in_buffer[96]<<0)-(in_buffer[96]<<2)-(in_buffer[96]<<4)-(in_buffer[96]<<6)+(in_buffer[96]<<11)+(in_buffer[96]<<12))-(0+(in_buffer[97]<<1)+(in_buffer[97]<<7)+(in_buffer[97]<<8)+(in_buffer[97]<<12))-(0+(in_buffer[98]<<2)+(in_buffer[98]<<3)+(in_buffer[98]<<6)+(in_buffer[98]<<8))-(0+(in_buffer[99]<<0)+(in_buffer[99]<<6)+(in_buffer[99]<<9)+(in_buffer[99]<<12)+(in_buffer[99]<<13))-(0+(in_buffer[100]<<0)+(in_buffer[100]<<4)+(in_buffer[100]<<8)-(in_buffer[100]<<10)+(in_buffer[100]<<12)+(in_buffer[100]<<13))-(0+(in_buffer[101]<<0)+(in_buffer[101]<<3)+(in_buffer[101]<<7)+(in_buffer[101]<<12))-(0+(in_buffer[102]<<3)-(in_buffer[102]<<6)+(in_buffer[102]<<11))-(0+(in_buffer[103]<<0)+(in_buffer[103]<<6)+(in_buffer[103]<<7)+(in_buffer[103]<<11))+(0+(in_buffer[104]<<1)+(in_buffer[104]<<2)-(in_buffer[104]<<8)+(in_buffer[104]<<10)+(in_buffer[104]<<11))-(0+(in_buffer[105]<<1)+(in_buffer[105]<<3)+(in_buffer[105]<<7)+(in_buffer[105]<<10))+(0+(in_buffer[106]<<0)+(in_buffer[106]<<4)-(in_buffer[106]<<7)+(in_buffer[106]<<10))-(0-(in_buffer[107]<<1)-(in_buffer[107]<<3)+(in_buffer[107]<<6)+(in_buffer[107]<<12))-(0+(in_buffer[108]<<0)-(in_buffer[108]<<4)-(in_buffer[108]<<6)+(in_buffer[108]<<8)+(in_buffer[108]<<9)+(in_buffer[108]<<13))-(0+(in_buffer[109]<<0)+(in_buffer[109]<<2)+(in_buffer[109]<<3)-(in_buffer[109]<<7)+(in_buffer[109]<<10)+(in_buffer[109]<<12)+(in_buffer[109]<<13))-(0-(in_buffer[110]<<3)+(in_buffer[110]<<7)-(in_buffer[110]<<9)-(in_buffer[110]<<11)+(in_buffer[110]<<14))-(0+(in_buffer[111]<<5)+(in_buffer[111]<<6)+(in_buffer[111]<<9)+(in_buffer[111]<<11))+(0+(in_buffer[112]<<5)+(in_buffer[112]<<6)+(in_buffer[112]<<9)+(in_buffer[112]<<11))-(0+(in_buffer[113]<<1)+(in_buffer[113]<<7)+(in_buffer[113]<<8)+(in_buffer[113]<<12))+(0-(in_buffer[114]<<0)+(in_buffer[114]<<3)+(in_buffer[114]<<4)+(in_buffer[114]<<7)-(in_buffer[114]<<9)+(in_buffer[114]<<12))+(0+(in_buffer[115]<<0)+(in_buffer[115]<<1)-(in_buffer[115]<<8)+(in_buffer[115]<<12)+(in_buffer[115]<<13))+(0+(in_buffer[116]<<0)+(in_buffer[116]<<2)+(in_buffer[116]<<5)+(in_buffer[116]<<7)+(in_buffer[116]<<10)+(in_buffer[116]<<11))+(0+(in_buffer[117]<<0)-(in_buffer[117]<<3)+(in_buffer[117]<<8))-(0+(in_buffer[118]<<0)+(in_buffer[118]<<1)-(in_buffer[118]<<7)+(in_buffer[118]<<9)+(in_buffer[118]<<10))-(0-(in_buffer[119]<<0)+(in_buffer[119]<<4)+(in_buffer[119]<<5)+(in_buffer[119]<<8)+(in_buffer[119]<<12))-(0+(in_buffer[120]<<1)+(in_buffer[120]<<2)-(in_buffer[120]<<6)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<1)-(in_buffer[0]<<4)-(in_buffer[0]<<7)+(in_buffer[0]<<13))-(0-(in_buffer[1]<<2)-(in_buffer[1]<<4)+(in_buffer[1]<<7)+(in_buffer[1]<<13))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<1)-(in_buffer[2]<<7)+(in_buffer[2]<<9)+(in_buffer[2]<<10))+(0-(in_buffer[3]<<2)-(in_buffer[3]<<4)-(in_buffer[3]<<6)+(in_buffer[3]<<10)+(in_buffer[3]<<11))+(0-(in_buffer[4]<<1)+(in_buffer[4]<<4)-(in_buffer[4]<<6)+(in_buffer[4]<<8)+(in_buffer[4]<<9)+(in_buffer[4]<<12))+(0-(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<7)+(in_buffer[5]<<9)+(in_buffer[5]<<12))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<6)+(in_buffer[6]<<7)+(in_buffer[6]<<13))+(0-(in_buffer[7]<<1)+(in_buffer[7]<<6)+(in_buffer[7]<<8)+(in_buffer[7]<<9))+(0-(in_buffer[8]<<0)-(in_buffer[8]<<2)-(in_buffer[8]<<4)+(in_buffer[8]<<8)+(in_buffer[8]<<9))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<1)-(in_buffer[9]<<7)+(in_buffer[9]<<9)+(in_buffer[9]<<10))+(0+(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<10)+(in_buffer[10]<<13))+(0-(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<4)+(in_buffer[11]<<7)+(in_buffer[11]<<9)+(in_buffer[11]<<11)+(in_buffer[11]<<12))+(0-(in_buffer[12]<<1)+(in_buffer[12]<<4)-(in_buffer[12]<<7)+(in_buffer[12]<<11)+(in_buffer[12]<<13))+(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<6)-(in_buffer[13]<<8)+(in_buffer[13]<<11)+(in_buffer[13]<<13))-(0+(in_buffer[14]<<1)-(in_buffer[14]<<4)+(in_buffer[14]<<9))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<2)-(in_buffer[15]<<4)-(in_buffer[15]<<7)+(in_buffer[15]<<11))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<1)-(in_buffer[16]<<7)+(in_buffer[16]<<9)+(in_buffer[16]<<10))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4)+(in_buffer[17]<<6))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<3)+(in_buffer[18]<<7)+(in_buffer[18]<<10))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<5)+(in_buffer[19]<<8)+(in_buffer[19]<<9)+(in_buffer[19]<<12))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<3)-(in_buffer[20]<<9)+(in_buffer[20]<<12)+(in_buffer[20]<<13))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<4)-(in_buffer[21]<<7)+(in_buffer[21]<<10))+(0+(in_buffer[22]<<2)+(in_buffer[22]<<4)+(in_buffer[22]<<5)+(in_buffer[22]<<11)+(in_buffer[22]<<13))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)-(in_buffer[23]<<8)+(in_buffer[23]<<11)+(in_buffer[23]<<12))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<5)-(in_buffer[24]<<9)+(in_buffer[24]<<13))+(0+(in_buffer[25]<<2)+(in_buffer[25]<<6)-(in_buffer[25]<<9)+(in_buffer[25]<<12))-(0+(in_buffer[26]<<1)+(in_buffer[26]<<3)-(in_buffer[26]<<5)-(in_buffer[26]<<8)+(in_buffer[26]<<12))-(0+(in_buffer[27]<<2)+(in_buffer[27]<<6)-(in_buffer[27]<<9)+(in_buffer[27]<<12))-(0-(in_buffer[28]<<1)-(in_buffer[28]<<4)+(in_buffer[28]<<7)+(in_buffer[28]<<11))+(0+(in_buffer[29]<<1)+(in_buffer[29]<<3)+(in_buffer[29]<<7)+(in_buffer[29]<<10))+(0+(in_buffer[30]<<0)+(in_buffer[30]<<2)+(in_buffer[30]<<5)+(in_buffer[30]<<7)+(in_buffer[30]<<10)+(in_buffer[30]<<11))+(0-(in_buffer[31]<<3)+(in_buffer[31]<<8)+(in_buffer[31]<<10)+(in_buffer[31]<<11))+(0+(in_buffer[32]<<1)+(in_buffer[32]<<2)-(in_buffer[32]<<8)+(in_buffer[32]<<10)+(in_buffer[32]<<11))+(0-(in_buffer[33]<<1)-(in_buffer[33]<<3)+(in_buffer[33]<<8)+(in_buffer[33]<<10)+(in_buffer[33]<<13))+(0+(in_buffer[34]<<2)+(in_buffer[34]<<4)+(in_buffer[34]<<8)+(in_buffer[34]<<11))+(0+(in_buffer[35]<<0)+(in_buffer[35]<<3)+(in_buffer[35]<<4)+(in_buffer[35]<<13))+(0+(in_buffer[36]<<1)-(in_buffer[36]<<3)-(in_buffer[36]<<5)+(in_buffer[36]<<8)+(in_buffer[36]<<11)+(in_buffer[36]<<13))+(0-(in_buffer[37]<<1)-(in_buffer[37]<<3)+(in_buffer[37]<<6)+(in_buffer[37]<<12))-(0+(in_buffer[38]<<0)+(in_buffer[38]<<2)-(in_buffer[38]<<4)-(in_buffer[38]<<7)+(in_buffer[38]<<11))+(0-(in_buffer[39]<<0)-(in_buffer[39]<<2)+(in_buffer[39]<<5)+(in_buffer[39]<<11))+(0+(in_buffer[40]<<1)+(in_buffer[40]<<2)-(in_buffer[40]<<5)-(in_buffer[40]<<7)-(in_buffer[40]<<9)+(in_buffer[40]<<11)+(in_buffer[40]<<12))+(0-(in_buffer[41]<<0)-(in_buffer[41]<<2)+(in_buffer[41]<<7)+(in_buffer[41]<<9)+(in_buffer[41]<<12))-(0-(in_buffer[42]<<1)+(in_buffer[42]<<6)+(in_buffer[42]<<8)+(in_buffer[42]<<9))+(0+(in_buffer[43]<<0)+(in_buffer[43]<<2)+(in_buffer[43]<<6)+(in_buffer[43]<<9))+(0+(in_buffer[44]<<1)+(in_buffer[44]<<4)+(in_buffer[44]<<8)+(in_buffer[44]<<13))-(0+(in_buffer[45]<<0)-(in_buffer[45]<<2)-(in_buffer[45]<<4)+(in_buffer[45]<<7)+(in_buffer[45]<<10)+(in_buffer[45]<<12))-(0+(in_buffer[46]<<0)-(in_buffer[46]<<3)+(in_buffer[46]<<8))+(0-(in_buffer[47]<<1)+(in_buffer[47]<<4)-(in_buffer[47]<<6)+(in_buffer[47]<<8)+(in_buffer[47]<<9)+(in_buffer[47]<<12))+(0+(in_buffer[48]<<0)+(in_buffer[48]<<3)+(in_buffer[48]<<7)+(in_buffer[48]<<12))-(0+(in_buffer[49]<<2)-(in_buffer[49]<<5)+(in_buffer[49]<<10))+(0+(in_buffer[50]<<0)+(in_buffer[50]<<6)+(in_buffer[50]<<7)+(in_buffer[50]<<11))+(0+(in_buffer[51]<<0)+(in_buffer[51]<<2)-(in_buffer[51]<<8)+(in_buffer[51]<<11)+(in_buffer[51]<<12))+(0+(in_buffer[52]<<1)-(in_buffer[52]<<5)-(in_buffer[52]<<10)+(in_buffer[52]<<13))+(0+(in_buffer[53]<<1)-(in_buffer[53]<<4)+(in_buffer[53]<<9))-(0+(in_buffer[54]<<0)+(in_buffer[54]<<6)+(in_buffer[54]<<7)+(in_buffer[54]<<11))-(0+(in_buffer[55]<<0)+(in_buffer[55]<<2)+(in_buffer[55]<<3)+(in_buffer[55]<<9)+(in_buffer[55]<<11))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<5)+(in_buffer[56]<<7)+(in_buffer[56]<<10)+(in_buffer[56]<<11))-(0+(in_buffer[57]<<4)-(in_buffer[57]<<7)+(in_buffer[57]<<12))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<3)+(in_buffer[58]<<5)+(in_buffer[58]<<9)+(in_buffer[58]<<10))+(0+(in_buffer[59]<<0)+(in_buffer[59]<<6)+(in_buffer[59]<<7)+(in_buffer[59]<<11))-(0-(in_buffer[60]<<1)-(in_buffer[60]<<3)-(in_buffer[60]<<5)+(in_buffer[60]<<9)+(in_buffer[60]<<10))+(0+(in_buffer[61]<<2)+(in_buffer[61]<<6)-(in_buffer[61]<<9)+(in_buffer[61]<<12))+(0-(in_buffer[62]<<0)+(in_buffer[62]<<3)-(in_buffer[62]<<5)+(in_buffer[62]<<7)+(in_buffer[62]<<8)+(in_buffer[62]<<11))+(0+(in_buffer[63]<<0)+(in_buffer[63]<<1)-(in_buffer[63]<<4)-(in_buffer[63]<<6)-(in_buffer[63]<<8)+(in_buffer[63]<<10)+(in_buffer[63]<<11))-(0-(in_buffer[64]<<1)-(in_buffer[64]<<3)-(in_buffer[64]<<5)+(in_buffer[64]<<9)+(in_buffer[64]<<10))-(0-(in_buffer[66]<<0)+(in_buffer[66]<<4)-(in_buffer[66]<<7)-(in_buffer[66]<<10)+(in_buffer[66]<<13))+(0+(in_buffer[67]<<0)-(in_buffer[67]<<2)+(in_buffer[67]<<6)-(in_buffer[67]<<8)+(in_buffer[67]<<12))-(0-(in_buffer[68]<<1)+(in_buffer[68]<<5)-(in_buffer[68]<<7)-(in_buffer[68]<<9)+(in_buffer[68]<<12))-(0-(in_buffer[69]<<2)-(in_buffer[69]<<4)-(in_buffer[69]<<6)+(in_buffer[69]<<10)+(in_buffer[69]<<11))+(0+(in_buffer[70]<<1)+(in_buffer[70]<<4)+(in_buffer[70]<<6)+(in_buffer[70]<<10)+(in_buffer[70]<<11))-(0+(in_buffer[71]<<0)+(in_buffer[71]<<2)+(in_buffer[71]<<6)+(in_buffer[71]<<9))+(0+(in_buffer[72]<<1)-(in_buffer[72]<<3)-(in_buffer[72]<<6)+(in_buffer[72]<<9)+(in_buffer[72]<<11))-(0+(in_buffer[73]<<1)-(in_buffer[73]<<3)-(in_buffer[73]<<6)+(in_buffer[73]<<9)+(in_buffer[73]<<11))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<3)+(in_buffer[74]<<8))+(0+(in_buffer[75]<<0)+(in_buffer[75]<<2)+(in_buffer[75]<<6)+(in_buffer[75]<<9))+(0-(in_buffer[76]<<0)-(in_buffer[76]<<2)-(in_buffer[76]<<4)+(in_buffer[76]<<8)+(in_buffer[76]<<9))-(0+(in_buffer[77]<<2)+(in_buffer[77]<<4)+(in_buffer[77]<<8)+(in_buffer[77]<<11))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)-(in_buffer[78]<<4)+(in_buffer[78]<<8)+(in_buffer[78]<<9))-(0+(in_buffer[79]<<2)+(in_buffer[79]<<4)-(in_buffer[79]<<6)-(in_buffer[79]<<9)+(in_buffer[79]<<13))-(0+(in_buffer[80]<<0)+(in_buffer[80]<<2)+(in_buffer[80]<<5)+(in_buffer[80]<<7)+(in_buffer[80]<<10)+(in_buffer[80]<<11))+(0+(in_buffer[81]<<1)-(in_buffer[81]<<3)-(in_buffer[81]<<6)+(in_buffer[81]<<9)+(in_buffer[81]<<11))-(0+(in_buffer[82]<<3)+(in_buffer[82]<<4)+(in_buffer[82]<<7)+(in_buffer[82]<<9))+(0+(in_buffer[83]<<0)+(in_buffer[83]<<2)-(in_buffer[83]<<4)-(in_buffer[83]<<7)+(in_buffer[83]<<11))-(0-(in_buffer[84]<<0)+(in_buffer[84]<<2)+(in_buffer[84]<<3)+(in_buffer[84]<<6)+(in_buffer[84]<<8)+(in_buffer[84]<<10)+(in_buffer[84]<<11))-(0-(in_buffer[85]<<1)+(in_buffer[85]<<6)+(in_buffer[85]<<8)+(in_buffer[85]<<9))+(0+(in_buffer[86]<<0)-(in_buffer[86]<<2)-(in_buffer[86]<<5)+(in_buffer[86]<<8)+(in_buffer[86]<<10))+(0+(in_buffer[87]<<1)-(in_buffer[87]<<4)+(in_buffer[87]<<9))+(0+(in_buffer[88]<<1)-(in_buffer[88]<<4)+(in_buffer[88]<<9))+(0+(in_buffer[89]<<1)+(in_buffer[89]<<5)-(in_buffer[89]<<8)+(in_buffer[89]<<11))-(0-(in_buffer[90]<<0)-(in_buffer[90]<<3)+(in_buffer[90]<<8)+(in_buffer[90]<<11)+(in_buffer[90]<<12))-(0-(in_buffer[91]<<0)+(in_buffer[91]<<4)+(in_buffer[91]<<5)+(in_buffer[91]<<8)+(in_buffer[91]<<12))+(0+(in_buffer[92]<<0)+(in_buffer[92]<<1)-(in_buffer[92]<<5)+(in_buffer[92]<<12))+(0+(in_buffer[93]<<3)-(in_buffer[93]<<6)+(in_buffer[93]<<11))-(0-(in_buffer[94]<<0)+(in_buffer[94]<<5)+(in_buffer[94]<<7)+(in_buffer[94]<<8))-(0-(in_buffer[95]<<0)-(in_buffer[95]<<3)+(in_buffer[95]<<6)+(in_buffer[95]<<10))-(0+(in_buffer[96]<<0)+(in_buffer[96]<<1)+(in_buffer[96]<<4)+(in_buffer[96]<<6))-(0+(in_buffer[97]<<0)+(in_buffer[97]<<2)-(in_buffer[97]<<4)-(in_buffer[97]<<7)+(in_buffer[97]<<11))-(0+(in_buffer[98]<<1)-(in_buffer[98]<<3)-(in_buffer[98]<<6)+(in_buffer[98]<<9)+(in_buffer[98]<<11))+(0-(in_buffer[99]<<0)+(in_buffer[99]<<3)-(in_buffer[99]<<5)+(in_buffer[99]<<7)+(in_buffer[99]<<8)+(in_buffer[99]<<11))+(0-(in_buffer[100]<<0)+(in_buffer[100]<<4)-(in_buffer[100]<<6)-(in_buffer[100]<<8)+(in_buffer[100]<<11))-(0+(in_buffer[101]<<0)+(in_buffer[101]<<2)+(in_buffer[101]<<3)+(in_buffer[101]<<9)+(in_buffer[101]<<11))-(0+(in_buffer[102]<<0)-(in_buffer[102]<<3)-(in_buffer[102]<<6)-(in_buffer[102]<<9)+(in_buffer[102]<<11)+(in_buffer[102]<<12))+(0+(in_buffer[103]<<0)+(in_buffer[103]<<4)-(in_buffer[103]<<7)+(in_buffer[103]<<10))+(0-(in_buffer[104]<<1)-(in_buffer[104]<<3)-(in_buffer[104]<<5)+(in_buffer[104]<<9)+(in_buffer[104]<<10))+(0+(in_buffer[105]<<0)-(in_buffer[105]<<2)-(in_buffer[105]<<5)+(in_buffer[105]<<8)+(in_buffer[105]<<10))-(0+(in_buffer[106]<<0)+(in_buffer[106]<<2)+(in_buffer[106]<<3)+(in_buffer[106]<<9)+(in_buffer[106]<<11))-(0+(in_buffer[107]<<0)+(in_buffer[107]<<1)+(in_buffer[107]<<4)+(in_buffer[107]<<8)+(in_buffer[107]<<10)+(in_buffer[107]<<12))-(0-(in_buffer[108]<<0)+(in_buffer[108]<<10)+(in_buffer[108]<<11))-(0+(in_buffer[109]<<4)-(in_buffer[109]<<7)+(in_buffer[109]<<12))+(0-(in_buffer[110]<<1)-(in_buffer[110]<<3)-(in_buffer[110]<<5)+(in_buffer[110]<<9)+(in_buffer[110]<<10))-(0+(in_buffer[111]<<5)+(in_buffer[111]<<6)+(in_buffer[111]<<9)+(in_buffer[111]<<11))+(0+(in_buffer[112]<<1)+(in_buffer[112]<<2)+(in_buffer[112]<<5)+(in_buffer[112]<<7))-(0+(in_buffer[113]<<1)-(in_buffer[113]<<5)-(in_buffer[113]<<10)+(in_buffer[113]<<13))-(0+(in_buffer[114]<<0)+(in_buffer[114]<<1)-(in_buffer[114]<<7)+(in_buffer[114]<<9)+(in_buffer[114]<<10))+(0+(in_buffer[115]<<0)+(in_buffer[115]<<3)+(in_buffer[115]<<7)+(in_buffer[115]<<12))+(0+(in_buffer[116]<<0)-(in_buffer[116]<<2)+(in_buffer[116]<<6)-(in_buffer[116]<<8)+(in_buffer[116]<<12))-(0+(in_buffer[117]<<2)+(in_buffer[117]<<4)+(in_buffer[117]<<8)+(in_buffer[117]<<11))-(0-(in_buffer[118]<<3)+(in_buffer[118]<<8)+(in_buffer[118]<<10)+(in_buffer[118]<<11))-(0+(in_buffer[119]<<3)-(in_buffer[119]<<6)+(in_buffer[119]<<11))-(0+(in_buffer[120]<<1)+(in_buffer[120]<<4)+(in_buffer[120]<<6)+(in_buffer[120]<<10)+(in_buffer[120]<<11));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0-(0+(in_buffer[0]<<2)+(in_buffer[0]<<3)-(in_buffer[0]<<6)-(in_buffer[0]<<8)-(in_buffer[0]<<10)+(in_buffer[0]<<12)+(in_buffer[0]<<13))+(0-(in_buffer[1]<<1)+(in_buffer[1]<<4)-(in_buffer[1]<<7)+(in_buffer[1]<<11)+(in_buffer[1]<<13))+(0-(in_buffer[2]<<0)-(in_buffer[2]<<2)+(in_buffer[2]<<7)+(in_buffer[2]<<9)+(in_buffer[2]<<12))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<2)-(in_buffer[3]<<8)+(in_buffer[3]<<10)+(in_buffer[3]<<11))-(0-(in_buffer[4]<<0)-(in_buffer[4]<<2)+(in_buffer[4]<<7)+(in_buffer[4]<<9)+(in_buffer[4]<<12))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<4)-(in_buffer[5]<<7)+(in_buffer[5]<<10))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<6)+(in_buffer[6]<<7)+(in_buffer[6]<<11))-(0-(in_buffer[7]<<1)-(in_buffer[7]<<4)+(in_buffer[7]<<7)+(in_buffer[7]<<11))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<3)-(in_buffer[8]<<5)-(in_buffer[8]<<8)-(in_buffer[8]<<10)+(in_buffer[8]<<13))+(0-(in_buffer[9]<<4)-(in_buffer[9]<<7)+(in_buffer[9]<<10)+(in_buffer[9]<<14))+(0-(in_buffer[10]<<4)-(in_buffer[10]<<7)+(in_buffer[10]<<10)+(in_buffer[10]<<14))-(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<5)+(in_buffer[11]<<11))-(0+(in_buffer[12]<<3)+(in_buffer[12]<<5)+(in_buffer[12]<<9)+(in_buffer[12]<<12))-(0-(in_buffer[13]<<1)-(in_buffer[13]<<3)-(in_buffer[13]<<5)+(in_buffer[13]<<9)+(in_buffer[13]<<10))+(0+(in_buffer[14]<<3)+(in_buffer[14]<<4)+(in_buffer[14]<<7)+(in_buffer[14]<<9))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<4)-(in_buffer[15]<<6)-(in_buffer[15]<<8)+(in_buffer[15]<<11))+(0-(in_buffer[16]<<1)+(in_buffer[16]<<5)-(in_buffer[16]<<7)-(in_buffer[16]<<9)+(in_buffer[16]<<12))+(0+(in_buffer[17]<<1)+(in_buffer[17]<<3)+(in_buffer[17]<<7)+(in_buffer[17]<<10))+(0+(in_buffer[18]<<1)-(in_buffer[18]<<4)+(in_buffer[18]<<9))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<10)+(in_buffer[19]<<11))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<5)+(in_buffer[20]<<7)+(in_buffer[20]<<10)+(in_buffer[20]<<11))+(0+(in_buffer[21]<<0)-(in_buffer[21]<<3)-(in_buffer[21]<<5)+(in_buffer[21]<<8)+(in_buffer[21]<<10)+(in_buffer[21]<<12)+(in_buffer[21]<<13))+(0+(in_buffer[22]<<2)-(in_buffer[22]<<4)-(in_buffer[22]<<7)+(in_buffer[22]<<10)+(in_buffer[22]<<12))-(0+(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<7)+(in_buffer[23]<<11)+(in_buffer[23]<<12))-(0+(in_buffer[24]<<3)-(in_buffer[24]<<6)+(in_buffer[24]<<11))-(0+(in_buffer[25]<<0)+(in_buffer[25]<<2)-(in_buffer[25]<<8)+(in_buffer[25]<<11)+(in_buffer[25]<<12))+(0-(in_buffer[26]<<1)-(in_buffer[26]<<3)+(in_buffer[26]<<6)+(in_buffer[26]<<12))+(0+(in_buffer[27]<<1)+(in_buffer[27]<<7)+(in_buffer[27]<<8)+(in_buffer[27]<<12))+(0+(in_buffer[28]<<1)+(in_buffer[28]<<4)+(in_buffer[28]<<6)+(in_buffer[28]<<10)+(in_buffer[28]<<11))-(0-(in_buffer[29]<<1)-(in_buffer[29]<<4)+(in_buffer[29]<<7)+(in_buffer[29]<<11))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<1)+(in_buffer[31]<<4)+(in_buffer[31]<<6))+(0-(in_buffer[32]<<0)+(in_buffer[32]<<2)+(in_buffer[32]<<3)+(in_buffer[32]<<9)+(in_buffer[32]<<13))+(0+(in_buffer[33]<<0)+(in_buffer[33]<<2)-(in_buffer[33]<<4)-(in_buffer[33]<<7)+(in_buffer[33]<<11))-(0+(in_buffer[34]<<1)+(in_buffer[34]<<7)+(in_buffer[34]<<8)+(in_buffer[34]<<12))-(0-(in_buffer[35]<<1)+(in_buffer[35]<<5)-(in_buffer[35]<<7)-(in_buffer[35]<<9)+(in_buffer[35]<<12))-(0+(in_buffer[36]<<2)+(in_buffer[36]<<4)+(in_buffer[36]<<5)+(in_buffer[36]<<11)+(in_buffer[36]<<13))-(0-(in_buffer[37]<<0)+(in_buffer[37]<<3)-(in_buffer[37]<<5)+(in_buffer[37]<<7)+(in_buffer[37]<<8)+(in_buffer[37]<<11))+(0-(in_buffer[38]<<1)+(in_buffer[38]<<5)-(in_buffer[38]<<7)-(in_buffer[38]<<9)+(in_buffer[38]<<12))+(0+(in_buffer[39]<<0)+(in_buffer[39]<<3)+(in_buffer[39]<<5)+(in_buffer[39]<<9)+(in_buffer[39]<<10))-(0+(in_buffer[40]<<2)+(in_buffer[40]<<6)-(in_buffer[40]<<9)+(in_buffer[40]<<12))-(0-(in_buffer[41]<<0)+(in_buffer[41]<<4)-(in_buffer[41]<<6)-(in_buffer[41]<<8)+(in_buffer[41]<<11))+(0-(in_buffer[42]<<0)+(in_buffer[42]<<3)-(in_buffer[42]<<6)+(in_buffer[42]<<10)+(in_buffer[42]<<12))-(0-(in_buffer[43]<<1)-(in_buffer[43]<<4)+(in_buffer[43]<<7)+(in_buffer[43]<<11))-(0+(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<10)+(in_buffer[44]<<13))-(0+(in_buffer[45]<<2)+(in_buffer[45]<<4)+(in_buffer[45]<<8)+(in_buffer[45]<<11))-(0+(in_buffer[46]<<1)-(in_buffer[46]<<3)-(in_buffer[46]<<6)+(in_buffer[46]<<9)+(in_buffer[46]<<11))-(0-(in_buffer[47]<<0)+(in_buffer[47]<<3)-(in_buffer[47]<<6)+(in_buffer[47]<<10)+(in_buffer[47]<<12))-(0-(in_buffer[48]<<1)-(in_buffer[48]<<4)+(in_buffer[48]<<7)+(in_buffer[48]<<11))+(0+(in_buffer[49]<<0)-(in_buffer[49]<<3)-(in_buffer[49]<<5)-(in_buffer[49]<<7)+(in_buffer[49]<<10)+(in_buffer[49]<<11))-(0-(in_buffer[50]<<0)+(in_buffer[50]<<5)+(in_buffer[50]<<7)+(in_buffer[50]<<8))+(0+(in_buffer[51]<<0)-(in_buffer[51]<<3)+(in_buffer[51]<<8))+(0+(in_buffer[52]<<2)+(in_buffer[52]<<3)+(in_buffer[52]<<6)+(in_buffer[52]<<8))+(0-(in_buffer[53]<<1)+(in_buffer[53]<<3)+(in_buffer[53]<<4)+(in_buffer[53]<<7)+(in_buffer[53]<<9)+(in_buffer[53]<<11)+(in_buffer[53]<<12))-(0+(in_buffer[54]<<0)+(in_buffer[54]<<1)+(in_buffer[54]<<4)+(in_buffer[54]<<8)+(in_buffer[54]<<10)+(in_buffer[54]<<12))+(0+(in_buffer[55]<<3)-(in_buffer[55]<<6)+(in_buffer[55]<<11))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<1)+(in_buffer[56]<<4)+(in_buffer[56]<<6))-(0+(in_buffer[57]<<0)+(in_buffer[57]<<3)+(in_buffer[57]<<5)+(in_buffer[57]<<9)+(in_buffer[57]<<10))-(0+(in_buffer[58]<<2)+(in_buffer[58]<<4)+(in_buffer[58]<<8)+(in_buffer[58]<<11))-(0+(in_buffer[59]<<0)+(in_buffer[59]<<3)+(in_buffer[59]<<5)+(in_buffer[59]<<9)+(in_buffer[59]<<10))+(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)-(in_buffer[60]<<5)+(in_buffer[60]<<12))+(0+(in_buffer[61]<<0)-(in_buffer[61]<<3)+(in_buffer[61]<<8))+(0+(in_buffer[62]<<5)+(in_buffer[62]<<6)+(in_buffer[62]<<9)+(in_buffer[62]<<11))+(0+(in_buffer[63]<<0)-(in_buffer[63]<<2)-(in_buffer[63]<<5)+(in_buffer[63]<<8)+(in_buffer[63]<<10))+(0-(in_buffer[64]<<0)+(in_buffer[64]<<4)+(in_buffer[64]<<5)+(in_buffer[64]<<8)+(in_buffer[64]<<12))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<3)+(in_buffer[65]<<6)+(in_buffer[65]<<10))+(0-(in_buffer[66]<<1)+(in_buffer[66]<<6)+(in_buffer[66]<<7)-(in_buffer[66]<<10)+(in_buffer[66]<<12)+(in_buffer[66]<<13))+(0+(in_buffer[67]<<0)+(in_buffer[67]<<4)+(in_buffer[67]<<6)+(in_buffer[67]<<11)+(in_buffer[67]<<12))-(0-(in_buffer[68]<<0)-(in_buffer[68]<<3)+(in_buffer[68]<<6)+(in_buffer[68]<<10))-(0-(in_buffer[69]<<0)+(in_buffer[69]<<5)+(in_buffer[69]<<7)+(in_buffer[69]<<8))-(0+(in_buffer[70]<<0)+(in_buffer[70]<<4)-(in_buffer[70]<<7)+(in_buffer[70]<<10))-(0-(in_buffer[71]<<0)+(in_buffer[71]<<5)+(in_buffer[71]<<7)+(in_buffer[71]<<8))-(0+(in_buffer[72]<<0)+(in_buffer[72]<<1)-(in_buffer[72]<<7)+(in_buffer[72]<<9)+(in_buffer[72]<<10))+(0+(in_buffer[73]<<1)+(in_buffer[73]<<5)-(in_buffer[73]<<8)+(in_buffer[73]<<11))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<2)-(in_buffer[74]<<5)+(in_buffer[74]<<8)+(in_buffer[74]<<10))+(0+(in_buffer[75]<<0)-(in_buffer[75]<<4)-(in_buffer[75]<<9)+(in_buffer[75]<<12))-(0+(in_buffer[76]<<0)+(in_buffer[76]<<1)+(in_buffer[76]<<4)+(in_buffer[76]<<6))-(0+(in_buffer[77]<<0)+(in_buffer[77]<<2)+(in_buffer[77]<<5)+(in_buffer[77]<<7)+(in_buffer[77]<<10)+(in_buffer[77]<<11))+(0+(in_buffer[78]<<1)+(in_buffer[78]<<3)+(in_buffer[78]<<6)+(in_buffer[78]<<8)+(in_buffer[78]<<11)+(in_buffer[78]<<12))+(0-(in_buffer[79]<<0)+(in_buffer[79]<<10)+(in_buffer[79]<<11))+(0+(in_buffer[80]<<2)-(in_buffer[80]<<4)-(in_buffer[80]<<7)+(in_buffer[80]<<10)+(in_buffer[80]<<12))-(0-(in_buffer[81]<<0)+(in_buffer[81]<<5)+(in_buffer[81]<<7)+(in_buffer[81]<<8))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)-(in_buffer[82]<<4)+(in_buffer[82]<<8)+(in_buffer[82]<<9))-(0+(in_buffer[83]<<0)+(in_buffer[83]<<2)-(in_buffer[83]<<4)-(in_buffer[83]<<7)+(in_buffer[83]<<11))+(0+(in_buffer[84]<<0)+(in_buffer[84]<<2)-(in_buffer[84]<<8)+(in_buffer[84]<<11)+(in_buffer[84]<<12))+(0+(in_buffer[85]<<4)-(in_buffer[85]<<7)+(in_buffer[85]<<12))+(0-(in_buffer[86]<<0)+(in_buffer[86]<<2)+(in_buffer[86]<<3)+(in_buffer[86]<<6)+(in_buffer[86]<<8)+(in_buffer[86]<<10)+(in_buffer[86]<<11))-(0+(in_buffer[87]<<1)+(in_buffer[87]<<7)+(in_buffer[87]<<8)+(in_buffer[87]<<12))-(0-(in_buffer[88]<<0)+(in_buffer[88]<<3)+(in_buffer[88]<<4)+(in_buffer[88]<<7)-(in_buffer[88]<<9)+(in_buffer[88]<<12))+(0+(in_buffer[89]<<0)+(in_buffer[89]<<1)-(in_buffer[89]<<7)+(in_buffer[89]<<9)+(in_buffer[89]<<10))+(0-(in_buffer[90]<<3)-(in_buffer[90]<<5)-(in_buffer[90]<<7)+(in_buffer[90]<<11)+(in_buffer[90]<<12))+(0+(in_buffer[91]<<0)+(in_buffer[91]<<2)-(in_buffer[91]<<5)+(in_buffer[91]<<7)+(in_buffer[91]<<8)+(in_buffer[91]<<13))-(0-(in_buffer[92]<<0)+(in_buffer[92]<<3)-(in_buffer[92]<<5)+(in_buffer[92]<<7)+(in_buffer[92]<<8)+(in_buffer[92]<<11))-(0+(in_buffer[93]<<2)+(in_buffer[93]<<4)+(in_buffer[93]<<8)+(in_buffer[93]<<11))-(0+(in_buffer[94]<<0)+(in_buffer[94]<<4)+(in_buffer[94]<<6)+(in_buffer[94]<<11)+(in_buffer[94]<<12))+(0-(in_buffer[95]<<0)+(in_buffer[95]<<10)+(in_buffer[95]<<11))+(0+(in_buffer[96]<<0)+(in_buffer[96]<<3)+(in_buffer[96]<<4)+(in_buffer[96]<<13))+(0-(in_buffer[97]<<0)+(in_buffer[97]<<3)-(in_buffer[97]<<6)+(in_buffer[97]<<10)+(in_buffer[97]<<12))+(0+(in_buffer[98]<<0)+(in_buffer[98]<<1)-(in_buffer[98]<<5)+(in_buffer[98]<<12))+(0-(in_buffer[99]<<0)+(in_buffer[99]<<2)+(in_buffer[99]<<3)+(in_buffer[99]<<6)+(in_buffer[99]<<8)+(in_buffer[99]<<10)+(in_buffer[99]<<11))+(0+(in_buffer[100]<<0)+(in_buffer[100]<<2)+(in_buffer[100]<<6)+(in_buffer[100]<<9))+(0-(in_buffer[101]<<0)-(in_buffer[101]<<3)+(in_buffer[101]<<8)+(in_buffer[101]<<11)+(in_buffer[101]<<12))+(0+(in_buffer[102]<<3)+(in_buffer[102]<<7)-(in_buffer[102]<<10)+(in_buffer[102]<<13))-(0-(in_buffer[103]<<1)+(in_buffer[103]<<6)+(in_buffer[103]<<8)+(in_buffer[103]<<9))-(0+(in_buffer[104]<<4)+(in_buffer[104]<<5)+(in_buffer[104]<<8)+(in_buffer[104]<<10))-(0+(in_buffer[105]<<0)+(in_buffer[105]<<2)+(in_buffer[105]<<4)-(in_buffer[105]<<6)+(in_buffer[105]<<9)+(in_buffer[105]<<12))+(0+(in_buffer[106]<<3)-(in_buffer[106]<<6)+(in_buffer[106]<<11))+(0+(in_buffer[107]<<4)+(in_buffer[107]<<6)+(in_buffer[107]<<10)+(in_buffer[107]<<13))+(0-(in_buffer[108]<<1)+(in_buffer[108]<<5)-(in_buffer[108]<<7)-(in_buffer[108]<<9)+(in_buffer[108]<<12))+(0-(in_buffer[109]<<1)+(in_buffer[109]<<11)+(in_buffer[109]<<12))+(0-(in_buffer[110]<<1)-(in_buffer[110]<<3)-(in_buffer[110]<<5)+(in_buffer[110]<<9)+(in_buffer[110]<<10))+(0+(in_buffer[111]<<4)-(in_buffer[111]<<7)+(in_buffer[111]<<12))+(0+(in_buffer[112]<<0)+(in_buffer[112]<<1)-(in_buffer[112]<<5)+(in_buffer[112]<<12))+(0-(in_buffer[113]<<0)+(in_buffer[113]<<5)+(in_buffer[113]<<6)-(in_buffer[113]<<9)+(in_buffer[113]<<11)+(in_buffer[113]<<12))+(0+(in_buffer[114]<<3)-(in_buffer[114]<<6)+(in_buffer[114]<<11))+(0+(in_buffer[115]<<1)+(in_buffer[115]<<3)+(in_buffer[115]<<7)+(in_buffer[115]<<10))-(0+(in_buffer[116]<<0)+(in_buffer[116]<<2)-(in_buffer[116]<<4)-(in_buffer[116]<<7)+(in_buffer[116]<<11))-(0-(in_buffer[117]<<0)+(in_buffer[117]<<3)-(in_buffer[117]<<5)+(in_buffer[117]<<7)+(in_buffer[117]<<8)+(in_buffer[117]<<11))+(0+(in_buffer[118]<<3)+(in_buffer[118]<<4)+(in_buffer[118]<<7)+(in_buffer[118]<<9))+(0+(in_buffer[119]<<5)+(in_buffer[119]<<6)+(in_buffer[119]<<9)+(in_buffer[119]<<11))+(0+(in_buffer[120]<<0)+(in_buffer[120]<<2)-(in_buffer[120]<<4)-(in_buffer[120]<<7)+(in_buffer[120]<<11));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0+(0+(in_buffer[0]<<4)+(in_buffer[0]<<5)+(in_buffer[0]<<8)+(in_buffer[0]<<10))+(0+(in_buffer[1]<<0)-(in_buffer[1]<<2)+(in_buffer[1]<<6)+(in_buffer[1]<<9)+(in_buffer[1]<<13)+(in_buffer[1]<<14))+(0-(in_buffer[2]<<0)+(in_buffer[2]<<3)-(in_buffer[2]<<6)+(in_buffer[2]<<10)+(in_buffer[2]<<12))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<4)+(in_buffer[3]<<6)+(in_buffer[3]<<10)+(in_buffer[3]<<11))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<4)+(in_buffer[4]<<6)+(in_buffer[4]<<11)+(in_buffer[4]<<12))+(0+(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<5)+(in_buffer[5]<<9)+(in_buffer[5]<<10))+(0+(in_buffer[6]<<1)+(in_buffer[6]<<2)-(in_buffer[6]<<8)+(in_buffer[6]<<10)+(in_buffer[6]<<11))+(0-(in_buffer[7]<<1)-(in_buffer[7]<<3)-(in_buffer[7]<<5)+(in_buffer[7]<<9)+(in_buffer[7]<<10))-(0+(in_buffer[8]<<4)-(in_buffer[8]<<7)+(in_buffer[8]<<12))+(0-(in_buffer[9]<<2)+(in_buffer[9]<<7)+(in_buffer[9]<<9)+(in_buffer[9]<<10))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)-(in_buffer[10]<<5)+(in_buffer[10]<<12))-(0-(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3)-(in_buffer[11]<<6)-(in_buffer[11]<<8)-(in_buffer[11]<<11)+(in_buffer[11]<<14))-(0+(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<6)-(in_buffer[12]<<8)+(in_buffer[12]<<12))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<1)-(in_buffer[13]<<4)-(in_buffer[13]<<7)+(in_buffer[13]<<13))-(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<6)-(in_buffer[14]<<8)+(in_buffer[14]<<12))-(0+(in_buffer[15]<<0)-(in_buffer[15]<<2)-(in_buffer[15]<<5)+(in_buffer[15]<<8)+(in_buffer[15]<<10))+(0+(in_buffer[16]<<1)+(in_buffer[16]<<2)+(in_buffer[16]<<5)+(in_buffer[16]<<7))-(0+(in_buffer[17]<<1)+(in_buffer[17]<<7)+(in_buffer[17]<<8)+(in_buffer[17]<<12))-(0+(in_buffer[18]<<4)+(in_buffer[18]<<6)+(in_buffer[18]<<10)+(in_buffer[18]<<13))-(0+(in_buffer[19]<<0)-(in_buffer[19]<<3)-(in_buffer[19]<<5)+(in_buffer[19]<<8)+(in_buffer[19]<<10)+(in_buffer[19]<<12)+(in_buffer[19]<<13))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<5)+(in_buffer[20]<<8)+(in_buffer[20]<<9)+(in_buffer[20]<<12))+(0-(in_buffer[21]<<0)-(in_buffer[21]<<4)+(in_buffer[21]<<9)+(in_buffer[21]<<10)+(in_buffer[21]<<13))-(0-(in_buffer[22]<<4)+(in_buffer[22]<<8)-(in_buffer[22]<<10)-(in_buffer[22]<<12)+(in_buffer[22]<<15))-(0+(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<9)+(in_buffer[23]<<14))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<1)-(in_buffer[24]<<5)+(in_buffer[24]<<12))+(0+(in_buffer[25]<<0)+(in_buffer[25]<<3)+(in_buffer[25]<<5)+(in_buffer[25]<<9)+(in_buffer[25]<<10))+(0+(in_buffer[26]<<0)-(in_buffer[26]<<4)-(in_buffer[26]<<9)+(in_buffer[26]<<12))+(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)+(in_buffer[27]<<7)+(in_buffer[27]<<9)+(in_buffer[27]<<12))-(0+(in_buffer[28]<<1)+(in_buffer[28]<<3)+(in_buffer[28]<<7)+(in_buffer[28]<<10))-(0-(in_buffer[29]<<1)+(in_buffer[29]<<5)-(in_buffer[29]<<7)-(in_buffer[29]<<9)+(in_buffer[29]<<12))-(0+(in_buffer[30]<<0)+(in_buffer[30]<<2)-(in_buffer[30]<<4)-(in_buffer[30]<<7)+(in_buffer[30]<<11))+(0+(in_buffer[31]<<4)-(in_buffer[31]<<7)+(in_buffer[31]<<12))+(0-(in_buffer[32]<<1)-(in_buffer[32]<<3)+(in_buffer[32]<<6)+(in_buffer[32]<<12))-(0-(in_buffer[33]<<0)+(in_buffer[33]<<3)+(in_buffer[33]<<8)+(in_buffer[33]<<10)+(in_buffer[33]<<13)+(in_buffer[33]<<15))-(0-(in_buffer[34]<<1)-(in_buffer[34]<<3)-(in_buffer[34]<<6)+(in_buffer[34]<<9)-(in_buffer[34]<<11)+(in_buffer[34]<<14))-(0+(in_buffer[35]<<3)+(in_buffer[35]<<5)+(in_buffer[35]<<9)+(in_buffer[35]<<12))-(0-(in_buffer[36]<<0)+(in_buffer[36]<<10)+(in_buffer[36]<<11))+(0-(in_buffer[37]<<0)+(in_buffer[37]<<2)+(in_buffer[37]<<3)+(in_buffer[37]<<6)+(in_buffer[37]<<8)+(in_buffer[37]<<10)+(in_buffer[37]<<11))+(0-(in_buffer[38]<<1)+(in_buffer[38]<<4)+(in_buffer[38]<<5)+(in_buffer[38]<<8)-(in_buffer[38]<<10)+(in_buffer[38]<<13))-(0+(in_buffer[40]<<0)+(in_buffer[40]<<6)+(in_buffer[40]<<7)+(in_buffer[40]<<11))-(0+(in_buffer[41]<<1)+(in_buffer[41]<<3)+(in_buffer[41]<<7)+(in_buffer[41]<<10))+(0+(in_buffer[42]<<0)-(in_buffer[42]<<3)+(in_buffer[42]<<8))-(0+(in_buffer[43]<<0)-(in_buffer[43]<<7)-(in_buffer[43]<<9)+(in_buffer[43]<<13))-(0-(in_buffer[44]<<1)-(in_buffer[44]<<3)+(in_buffer[44]<<5)+(in_buffer[44]<<6)+(in_buffer[44]<<9)+(in_buffer[44]<<15))-(0+(in_buffer[45]<<0)+(in_buffer[45]<<1)+(in_buffer[45]<<4)+(in_buffer[45]<<8)+(in_buffer[45]<<10)+(in_buffer[45]<<12))+(0-(in_buffer[46]<<1)-(in_buffer[46]<<4)+(in_buffer[46]<<7)+(in_buffer[46]<<11))+(0-(in_buffer[47]<<2)-(in_buffer[47]<<4)-(in_buffer[47]<<6)+(in_buffer[47]<<10)+(in_buffer[47]<<11))-(0+(in_buffer[48]<<0)+(in_buffer[48]<<1)-(in_buffer[48]<<7)+(in_buffer[48]<<9)+(in_buffer[48]<<10))+(0+(in_buffer[49]<<0)+(in_buffer[49]<<6)+(in_buffer[49]<<7)+(in_buffer[49]<<11))+(0+(in_buffer[50]<<0)-(in_buffer[50]<<2)+(in_buffer[50]<<6)-(in_buffer[50]<<8)+(in_buffer[50]<<12))+(0+(in_buffer[51]<<2)-(in_buffer[51]<<5)+(in_buffer[51]<<10))+(0+(in_buffer[52]<<0)+(in_buffer[52]<<1)+(in_buffer[52]<<4)+(in_buffer[52]<<6))-(0+(in_buffer[54]<<1)-(in_buffer[54]<<8)-(in_buffer[54]<<10)+(in_buffer[54]<<14))-(0+(in_buffer[55]<<0)-(in_buffer[55]<<3)+(in_buffer[55]<<8))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<3)+(in_buffer[56]<<5)+(in_buffer[56]<<9)+(in_buffer[56]<<10))+(0-(in_buffer[57]<<1)+(in_buffer[57]<<4)+(in_buffer[57]<<5)+(in_buffer[57]<<8)-(in_buffer[57]<<10)+(in_buffer[57]<<13))+(0-(in_buffer[58]<<2)-(in_buffer[58]<<5)+(in_buffer[58]<<8)+(in_buffer[58]<<12))-(0+(in_buffer[59]<<1)+(in_buffer[59]<<3)+(in_buffer[59]<<7)+(in_buffer[59]<<10))+(0+(in_buffer[60]<<0)-(in_buffer[60]<<3)+(in_buffer[60]<<8))+(0+(in_buffer[61]<<5)+(in_buffer[61]<<6)+(in_buffer[61]<<9)+(in_buffer[61]<<11))-(0-(in_buffer[62]<<0)+(in_buffer[62]<<5)+(in_buffer[62]<<7)+(in_buffer[62]<<8))+(0+(in_buffer[63]<<5)+(in_buffer[63]<<6)+(in_buffer[63]<<9)+(in_buffer[63]<<11))-(0+(in_buffer[64]<<0)-(in_buffer[64]<<3)-(in_buffer[64]<<6)-(in_buffer[64]<<9)+(in_buffer[64]<<11)+(in_buffer[64]<<12))-(0-(in_buffer[65]<<1)+(in_buffer[65]<<3)+(in_buffer[65]<<4)+(in_buffer[65]<<10)+(in_buffer[65]<<14))+(0-(in_buffer[66]<<4)+(in_buffer[66]<<9)+(in_buffer[66]<<11)+(in_buffer[66]<<12))-(0+(in_buffer[67]<<2)+(in_buffer[67]<<6)-(in_buffer[67]<<9)+(in_buffer[67]<<12))+(0-(in_buffer[68]<<0)-(in_buffer[68]<<2)+(in_buffer[68]<<7)+(in_buffer[68]<<9)+(in_buffer[68]<<12))+(0-(in_buffer[69]<<1)+(in_buffer[69]<<6)+(in_buffer[69]<<8)+(in_buffer[69]<<9))+(0-(in_buffer[70]<<0)+(in_buffer[70]<<3)-(in_buffer[70]<<5)+(in_buffer[70]<<7)+(in_buffer[70]<<8)+(in_buffer[70]<<11))-(0+(in_buffer[71]<<5)+(in_buffer[71]<<6)+(in_buffer[71]<<9)+(in_buffer[71]<<11))+(0+(in_buffer[72]<<0)+(in_buffer[72]<<2)+(in_buffer[72]<<3)+(in_buffer[72]<<9)+(in_buffer[72]<<11))+(0+(in_buffer[73]<<0)+(in_buffer[73]<<4)-(in_buffer[73]<<7)+(in_buffer[73]<<10))+(0-(in_buffer[74]<<3)+(in_buffer[74]<<8)+(in_buffer[74]<<10)+(in_buffer[74]<<11))-(0+(in_buffer[75]<<6)+(in_buffer[75]<<7)+(in_buffer[75]<<10)+(in_buffer[75]<<12))-(0+(in_buffer[76]<<1)+(in_buffer[76]<<2)+(in_buffer[76]<<5)+(in_buffer[76]<<7))+(0-(in_buffer[77]<<2)-(in_buffer[77]<<5)+(in_buffer[77]<<8)+(in_buffer[77]<<12))-(0+(in_buffer[78]<<1)-(in_buffer[78]<<4)+(in_buffer[78]<<9))+(0+(in_buffer[79]<<0)+(in_buffer[79]<<4)+(in_buffer[79]<<6)+(in_buffer[79]<<11)+(in_buffer[79]<<12))-(0+(in_buffer[80]<<0)-(in_buffer[80]<<3)+(in_buffer[80]<<8))+(0+(in_buffer[81]<<5)+(in_buffer[81]<<6)+(in_buffer[81]<<9)+(in_buffer[81]<<11))-(0+(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<5)+(in_buffer[82]<<7)+(in_buffer[82]<<8)+(in_buffer[82]<<11)+(in_buffer[82]<<12))+(0+(in_buffer[83]<<1)+(in_buffer[83]<<3)+(in_buffer[83]<<7)+(in_buffer[83]<<10))-(0+(in_buffer[84]<<0)+(in_buffer[84]<<2)-(in_buffer[84]<<4)-(in_buffer[84]<<7)+(in_buffer[84]<<11))+(0+(in_buffer[85]<<3)-(in_buffer[85]<<6)+(in_buffer[85]<<11))+(0+(in_buffer[86]<<0)-(in_buffer[86]<<3)+(in_buffer[86]<<8))+(0+(in_buffer[87]<<0)-(in_buffer[87]<<2)+(in_buffer[87]<<6)-(in_buffer[87]<<8)+(in_buffer[87]<<12))+(0+(in_buffer[88]<<5)+(in_buffer[88]<<6)+(in_buffer[88]<<9)+(in_buffer[88]<<11))-(0+(in_buffer[89]<<3)+(in_buffer[89]<<4)+(in_buffer[89]<<7)+(in_buffer[89]<<9))+(0+(in_buffer[90]<<1)-(in_buffer[90]<<3)-(in_buffer[90]<<6)+(in_buffer[90]<<9)+(in_buffer[90]<<11))-(0+(in_buffer[91]<<0)+(in_buffer[91]<<1)-(in_buffer[91]<<5)+(in_buffer[91]<<12))+(0+(in_buffer[92]<<4)-(in_buffer[92]<<7)+(in_buffer[92]<<12))-(0-(in_buffer[93]<<1)+(in_buffer[93]<<3)+(in_buffer[93]<<4)+(in_buffer[93]<<7)+(in_buffer[93]<<9)+(in_buffer[93]<<11)+(in_buffer[93]<<12))+(0-(in_buffer[94]<<1)+(in_buffer[94]<<5)-(in_buffer[94]<<7)-(in_buffer[94]<<9)+(in_buffer[94]<<12))-(0+(in_buffer[95]<<1)+(in_buffer[95]<<3)+(in_buffer[95]<<4)+(in_buffer[95]<<10)+(in_buffer[95]<<12))-(0+(in_buffer[96]<<1)+(in_buffer[96]<<5)-(in_buffer[96]<<8)+(in_buffer[96]<<11))-(0-(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<5)+(in_buffer[97]<<11))-(0-(in_buffer[98]<<0)+(in_buffer[98]<<5)+(in_buffer[98]<<7)+(in_buffer[98]<<8))-(0-(in_buffer[99]<<3)+(in_buffer[99]<<7)-(in_buffer[99]<<9)-(in_buffer[99]<<11)+(in_buffer[99]<<14))-(0+(in_buffer[100]<<0)-(in_buffer[100]<<2)+(in_buffer[100]<<10)+(in_buffer[100]<<13))+(0-(in_buffer[101]<<0)+(in_buffer[101]<<4)-(in_buffer[101]<<6)-(in_buffer[101]<<8)+(in_buffer[101]<<11))-(0+(in_buffer[102]<<0)+(in_buffer[102]<<1)-(in_buffer[102]<<5)+(in_buffer[102]<<12))+(0-(in_buffer[103]<<1)-(in_buffer[103]<<3)+(in_buffer[103]<<6)+(in_buffer[103]<<12))-(0-(in_buffer[104]<<0)+(in_buffer[104]<<3)-(in_buffer[104]<<6)+(in_buffer[104]<<10)+(in_buffer[104]<<12))+(0-(in_buffer[105]<<0)-(in_buffer[105]<<2)-(in_buffer[105]<<4)+(in_buffer[105]<<8)+(in_buffer[105]<<9))-(0-(in_buffer[106]<<0)+(in_buffer[106]<<5)+(in_buffer[106]<<6)-(in_buffer[106]<<9)+(in_buffer[106]<<11)+(in_buffer[106]<<12))+(0+(in_buffer[107]<<5)+(in_buffer[107]<<6)+(in_buffer[107]<<9)+(in_buffer[107]<<11))+(0-(in_buffer[108]<<1)-(in_buffer[108]<<3)-(in_buffer[108]<<5)+(in_buffer[108]<<9)+(in_buffer[108]<<10))-(0+(in_buffer[109]<<2)+(in_buffer[109]<<3)+(in_buffer[109]<<6)+(in_buffer[109]<<8))-(0+(in_buffer[110]<<1)-(in_buffer[110]<<5)-(in_buffer[110]<<10)+(in_buffer[110]<<13))-(0-(in_buffer[111]<<3)+(in_buffer[111]<<8)+(in_buffer[111]<<10)+(in_buffer[111]<<11))-(0+(in_buffer[112]<<0)+(in_buffer[112]<<6)+(in_buffer[112]<<7)+(in_buffer[112]<<11))-(0+(in_buffer[113]<<3)+(in_buffer[113]<<5)+(in_buffer[113]<<9)+(in_buffer[113]<<12))+(0-(in_buffer[114]<<2)-(in_buffer[114]<<4)-(in_buffer[114]<<6)+(in_buffer[114]<<10)+(in_buffer[114]<<11))-(0+(in_buffer[115]<<0)+(in_buffer[115]<<2)+(in_buffer[115]<<4)+(in_buffer[115]<<7)+(in_buffer[115]<<9)+(in_buffer[115]<<10)+(in_buffer[115]<<13))+(0+(in_buffer[116]<<0)+(in_buffer[116]<<1)+(in_buffer[116]<<4)+(in_buffer[116]<<8)+(in_buffer[116]<<10)+(in_buffer[116]<<12))+(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<5)+(in_buffer[118]<<11))+(0+(in_buffer[119]<<3)+(in_buffer[119]<<4)+(in_buffer[119]<<7)+(in_buffer[119]<<9))-(0-(in_buffer[120]<<1)+(in_buffer[120]<<4)+(in_buffer[120]<<5)+(in_buffer[120]<<8)-(in_buffer[120]<<10)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0+(0+(in_buffer[0]<<1)+(in_buffer[0]<<4)+(in_buffer[0]<<8)+(in_buffer[0]<<13))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<6)+(in_buffer[1]<<9))-(0+(in_buffer[2]<<0)-(in_buffer[2]<<4)-(in_buffer[2]<<9)+(in_buffer[2]<<12))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<4)+(in_buffer[3]<<6)+(in_buffer[3]<<10)+(in_buffer[3]<<11))+(0+(in_buffer[4]<<4)+(in_buffer[4]<<5)+(in_buffer[4]<<8)+(in_buffer[4]<<10))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<4)-(in_buffer[5]<<6)+(in_buffer[5]<<9)+(in_buffer[5]<<12))-(0-(in_buffer[6]<<2)-(in_buffer[6]<<4)-(in_buffer[6]<<6)+(in_buffer[6]<<10)+(in_buffer[6]<<11))-(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)-(in_buffer[7]<<4)-(in_buffer[7]<<6)+(in_buffer[7]<<11)+(in_buffer[7]<<12))-(0+(in_buffer[8]<<0)+(in_buffer[8]<<3)-(in_buffer[8]<<5)-(in_buffer[8]<<8)-(in_buffer[8]<<10)+(in_buffer[8]<<13))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<2)-(in_buffer[9]<<8)+(in_buffer[9]<<10)+(in_buffer[9]<<11))+(0-(in_buffer[10]<<0)+(in_buffer[10]<<5)+(in_buffer[10]<<7)+(in_buffer[10]<<8))-(0-(in_buffer[11]<<1)+(in_buffer[11]<<4)+(in_buffer[11]<<5)+(in_buffer[11]<<8)-(in_buffer[11]<<10)+(in_buffer[11]<<13))+(0+(in_buffer[12]<<0)-(in_buffer[12]<<2)-(in_buffer[12]<<4)+(in_buffer[12]<<7)+(in_buffer[12]<<10)+(in_buffer[12]<<12))-(0+(in_buffer[13]<<4)-(in_buffer[13]<<7)+(in_buffer[13]<<12))+(0-(in_buffer[14]<<1)-(in_buffer[14]<<3)+(in_buffer[14]<<6)+(in_buffer[14]<<12))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3)-(in_buffer[15]<<5)+(in_buffer[15]<<7)+(in_buffer[15]<<8)+(in_buffer[15]<<11))+(0+(in_buffer[16]<<0)+(in_buffer[16]<<5)+(in_buffer[16]<<8)+(in_buffer[16]<<9)+(in_buffer[16]<<12))-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)-(in_buffer[18]<<4)+(in_buffer[18]<<8)+(in_buffer[18]<<9))+(0-(in_buffer[19]<<1)+(in_buffer[19]<<6)+(in_buffer[19]<<8)+(in_buffer[19]<<9))+(0-(in_buffer[20]<<2)-(in_buffer[20]<<4)-(in_buffer[20]<<6)+(in_buffer[20]<<10)+(in_buffer[20]<<11))+(0+(in_buffer[21]<<4)+(in_buffer[21]<<5)+(in_buffer[21]<<8)+(in_buffer[21]<<10))-(0-(in_buffer[22]<<2)-(in_buffer[22]<<5)+(in_buffer[22]<<8)+(in_buffer[22]<<12))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<4)+(in_buffer[23]<<7)+(in_buffer[23]<<9)+(in_buffer[23]<<10)+(in_buffer[23]<<13))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<1)+(in_buffer[24]<<6)+(in_buffer[24]<<9)+(in_buffer[24]<<11)+(in_buffer[24]<<12))+(0+(in_buffer[25]<<0)+(in_buffer[25]<<4)-(in_buffer[25]<<7)+(in_buffer[25]<<10))+(0-(in_buffer[26]<<0)+(in_buffer[26]<<4)-(in_buffer[26]<<6)-(in_buffer[26]<<8)+(in_buffer[26]<<11))+(0-(in_buffer[27]<<0)+(in_buffer[27]<<5)+(in_buffer[27]<<7)+(in_buffer[27]<<8))-(0-(in_buffer[28]<<2)-(in_buffer[28]<<4)-(in_buffer[28]<<6)+(in_buffer[28]<<10)+(in_buffer[28]<<11))-(0-(in_buffer[29]<<3)+(in_buffer[29]<<8)+(in_buffer[29]<<10)+(in_buffer[29]<<11))+(0+(in_buffer[30]<<2)+(in_buffer[30]<<3)+(in_buffer[30]<<6)+(in_buffer[30]<<8))+(0-(in_buffer[31]<<1)-(in_buffer[31]<<3)-(in_buffer[31]<<5)+(in_buffer[31]<<9)+(in_buffer[31]<<10))-(0+(in_buffer[32]<<0)+(in_buffer[32]<<1)+(in_buffer[32]<<6)+(in_buffer[32]<<9)+(in_buffer[32]<<11)+(in_buffer[32]<<12))-(0+(in_buffer[33]<<0)+(in_buffer[33]<<4)+(in_buffer[33]<<6)+(in_buffer[33]<<11)+(in_buffer[33]<<12))+(0+(in_buffer[34]<<6)+(in_buffer[34]<<7)+(in_buffer[34]<<10)+(in_buffer[34]<<12))-(0+(in_buffer[35]<<0)+(in_buffer[35]<<2)+(in_buffer[35]<<6)+(in_buffer[35]<<9))+(0-(in_buffer[36]<<4)+(in_buffer[36]<<9)+(in_buffer[36]<<11)+(in_buffer[36]<<12))-(0+(in_buffer[37]<<2)+(in_buffer[37]<<4)+(in_buffer[37]<<8)+(in_buffer[37]<<11))+(0-(in_buffer[38]<<0)+(in_buffer[38]<<10)+(in_buffer[38]<<11))-(0-(in_buffer[39]<<1)-(in_buffer[39]<<4)+(in_buffer[39]<<7)+(in_buffer[39]<<11))+(0+(in_buffer[40]<<0)+(in_buffer[40]<<1)-(in_buffer[40]<<7)+(in_buffer[40]<<9)+(in_buffer[40]<<10))+(0+(in_buffer[41]<<0)+(in_buffer[41]<<2)-(in_buffer[41]<<8)+(in_buffer[41]<<11)+(in_buffer[41]<<12))-(0+(in_buffer[42]<<0)+(in_buffer[42]<<1)-(in_buffer[42]<<5)+(in_buffer[42]<<12))-(0-(in_buffer[43]<<0)+(in_buffer[43]<<3)+(in_buffer[43]<<4)+(in_buffer[43]<<7)-(in_buffer[43]<<9)+(in_buffer[43]<<12))-(0+(in_buffer[44]<<1)+(in_buffer[44]<<3)+(in_buffer[44]<<4)+(in_buffer[44]<<10)+(in_buffer[44]<<12))+(0+(in_buffer[45]<<0)-(in_buffer[45]<<3)-(in_buffer[45]<<5)-(in_buffer[45]<<7)+(in_buffer[45]<<10)+(in_buffer[45]<<11))+(0+(in_buffer[46]<<1)+(in_buffer[46]<<6)+(in_buffer[46]<<9)+(in_buffer[46]<<10)+(in_buffer[46]<<13))+(0-(in_buffer[47]<<0)+(in_buffer[47]<<6)+(in_buffer[47]<<7)+(in_buffer[47]<<13))-(0+(in_buffer[48]<<1)-(in_buffer[48]<<3)+(in_buffer[48]<<7)-(in_buffer[48]<<9)+(in_buffer[48]<<13))-(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)-(in_buffer[49]<<4)-(in_buffer[49]<<6)+(in_buffer[49]<<11)+(in_buffer[49]<<12))-(0-(in_buffer[50]<<3)+(in_buffer[50]<<8)+(in_buffer[50]<<10)+(in_buffer[50]<<11))+(0-(in_buffer[51]<<1)+(in_buffer[51]<<5)-(in_buffer[51]<<7)-(in_buffer[51]<<9)+(in_buffer[51]<<12))+(0+(in_buffer[52]<<0)+(in_buffer[52]<<5)+(in_buffer[52]<<8)+(in_buffer[52]<<9)+(in_buffer[52]<<12))-(0+(in_buffer[53]<<1)-(in_buffer[53]<<3)-(in_buffer[53]<<6)+(in_buffer[53]<<9)+(in_buffer[53]<<11))-(0+(in_buffer[54]<<1)+(in_buffer[54]<<4)+(in_buffer[54]<<6)+(in_buffer[54]<<10)+(in_buffer[54]<<11))-(0+(in_buffer[55]<<0)+(in_buffer[55]<<2)+(in_buffer[55]<<5)-(in_buffer[55]<<9)-(in_buffer[55]<<11)+(in_buffer[55]<<14))-(0+(in_buffer[56]<<1)+(in_buffer[56]<<2)-(in_buffer[56]<<6)+(in_buffer[56]<<13))+(0-(in_buffer[57]<<1)+(in_buffer[57]<<6)+(in_buffer[57]<<7)-(in_buffer[57]<<10)+(in_buffer[57]<<12)+(in_buffer[57]<<13))+(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)-(in_buffer[58]<<4)-(in_buffer[58]<<7)+(in_buffer[58]<<11))-(0-(in_buffer[59]<<0)-(in_buffer[59]<<2)+(in_buffer[59]<<5)+(in_buffer[59]<<11))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)-(in_buffer[60]<<4)-(in_buffer[60]<<6)-(in_buffer[60]<<8)+(in_buffer[60]<<10)+(in_buffer[60]<<11))-(0+(in_buffer[61]<<4)-(in_buffer[61]<<7)+(in_buffer[61]<<12))+(0-(in_buffer[62]<<2)+(in_buffer[62]<<7)+(in_buffer[62]<<9)+(in_buffer[62]<<10))+(0+(in_buffer[63]<<0)+(in_buffer[63]<<4)-(in_buffer[63]<<7)+(in_buffer[63]<<10))-(0+(in_buffer[64]<<5)+(in_buffer[64]<<6)+(in_buffer[64]<<9)+(in_buffer[64]<<11))-(0+(in_buffer[65]<<0)+(in_buffer[65]<<2)-(in_buffer[65]<<8)+(in_buffer[65]<<11)+(in_buffer[65]<<12))-(0+(in_buffer[66]<<1)-(in_buffer[66]<<3)+(in_buffer[66]<<7)-(in_buffer[66]<<9)+(in_buffer[66]<<13))-(0+(in_buffer[67]<<0)+(in_buffer[67]<<2)-(in_buffer[67]<<5)+(in_buffer[67]<<7)+(in_buffer[67]<<8)+(in_buffer[67]<<13))+(0-(in_buffer[68]<<0)+(in_buffer[68]<<3)-(in_buffer[68]<<5)+(in_buffer[68]<<8)+(in_buffer[68]<<9)+(in_buffer[68]<<12)+(in_buffer[68]<<13))+(0+(in_buffer[69]<<1)+(in_buffer[69]<<7)+(in_buffer[69]<<8)+(in_buffer[69]<<12))-(0+(in_buffer[70]<<1)+(in_buffer[70]<<3)+(in_buffer[70]<<7)+(in_buffer[70]<<10))+(0+(in_buffer[71]<<0)+(in_buffer[71]<<1)-(in_buffer[71]<<7)+(in_buffer[71]<<9)+(in_buffer[71]<<10))-(0-(in_buffer[72]<<0)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0-(in_buffer[73]<<2)-(in_buffer[73]<<4)-(in_buffer[73]<<6)+(in_buffer[73]<<10)+(in_buffer[73]<<11))+(0-(in_buffer[74]<<2)-(in_buffer[74]<<5)+(in_buffer[74]<<8)+(in_buffer[74]<<12))-(0+(in_buffer[75]<<0)-(in_buffer[75]<<3)-(in_buffer[75]<<5)-(in_buffer[75]<<7)+(in_buffer[75]<<10)+(in_buffer[75]<<11))-(0+(in_buffer[77]<<0)+(in_buffer[77]<<3)-(in_buffer[77]<<5)-(in_buffer[77]<<8)-(in_buffer[77]<<10)+(in_buffer[77]<<13))-(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<7)+(in_buffer[78]<<9)+(in_buffer[78]<<12))+(0+(in_buffer[79]<<0)-(in_buffer[79]<<2)+(in_buffer[79]<<4)+(in_buffer[79]<<5)+(in_buffer[79]<<8)+(in_buffer[79]<<11)+(in_buffer[79]<<13))+(0-(in_buffer[80]<<1)-(in_buffer[80]<<4)+(in_buffer[80]<<7)+(in_buffer[80]<<11))-(0+(in_buffer[81]<<3)+(in_buffer[81]<<4)+(in_buffer[81]<<7)+(in_buffer[81]<<9))+(0+(in_buffer[82]<<0)+(in_buffer[82]<<2)+(in_buffer[82]<<3)+(in_buffer[82]<<9)+(in_buffer[82]<<11))-(0+(in_buffer[83]<<1)+(in_buffer[83]<<3)+(in_buffer[83]<<4)+(in_buffer[83]<<10)+(in_buffer[83]<<12))-(0-(in_buffer[84]<<1)-(in_buffer[84]<<4)+(in_buffer[84]<<7)+(in_buffer[84]<<11))-(0+(in_buffer[85]<<1)+(in_buffer[85]<<2)+(in_buffer[85]<<5)+(in_buffer[85]<<7))+(0+(in_buffer[86]<<1)-(in_buffer[86]<<3)-(in_buffer[86]<<6)+(in_buffer[86]<<9)+(in_buffer[86]<<11))-(0+(in_buffer[87]<<1)-(in_buffer[87]<<3)-(in_buffer[87]<<6)+(in_buffer[87]<<9)+(in_buffer[87]<<11))-(0+(in_buffer[88]<<2)+(in_buffer[88]<<3)-(in_buffer[88]<<9)+(in_buffer[88]<<11)+(in_buffer[88]<<12))-(0+(in_buffer[89]<<0)+(in_buffer[89]<<3)+(in_buffer[89]<<5)+(in_buffer[89]<<9)+(in_buffer[89]<<10))+(0-(in_buffer[90]<<1)-(in_buffer[90]<<3)+(in_buffer[90]<<8)+(in_buffer[90]<<10)+(in_buffer[90]<<13))+(0+(in_buffer[91]<<1)+(in_buffer[91]<<4)+(in_buffer[91]<<6)+(in_buffer[91]<<10)+(in_buffer[91]<<11))-(0+(in_buffer[92]<<1)+(in_buffer[92]<<2)+(in_buffer[92]<<5)+(in_buffer[92]<<7))+(0+(in_buffer[93]<<1)+(in_buffer[93]<<4)+(in_buffer[93]<<6)+(in_buffer[93]<<10)+(in_buffer[93]<<11))-(0+(in_buffer[94]<<0)+(in_buffer[94]<<5)+(in_buffer[94]<<8)+(in_buffer[94]<<9)+(in_buffer[94]<<12))-(0+(in_buffer[95]<<2)+(in_buffer[95]<<5)+(in_buffer[95]<<7)+(in_buffer[95]<<11)+(in_buffer[95]<<12))+(0+(in_buffer[96]<<1)+(in_buffer[96]<<3)+(in_buffer[96]<<7)+(in_buffer[96]<<10))+(0+(in_buffer[97]<<1)+(in_buffer[97]<<3)+(in_buffer[97]<<7)+(in_buffer[97]<<10))-(0+(in_buffer[98]<<3)-(in_buffer[98]<<6)+(in_buffer[98]<<11))+(0-(in_buffer[99]<<0)-(in_buffer[99]<<2)-(in_buffer[99]<<4)+(in_buffer[99]<<8)+(in_buffer[99]<<9))-(0+(in_buffer[100]<<0)+(in_buffer[100]<<1)+(in_buffer[100]<<4)+(in_buffer[100]<<6))+(0+(in_buffer[101]<<2)-(in_buffer[101]<<5)+(in_buffer[101]<<10))+(0-(in_buffer[102]<<0)+(in_buffer[102]<<5)+(in_buffer[102]<<7)+(in_buffer[102]<<8))+(0+(in_buffer[103]<<0)+(in_buffer[103]<<2)+(in_buffer[103]<<6)+(in_buffer[103]<<9))+(0+(in_buffer[104]<<0)+(in_buffer[104]<<1)-(in_buffer[104]<<4)-(in_buffer[104]<<6)-(in_buffer[104]<<8)+(in_buffer[104]<<10)+(in_buffer[104]<<11))+(0-(in_buffer[105]<<0)+(in_buffer[105]<<4)-(in_buffer[105]<<6)-(in_buffer[105]<<8)+(in_buffer[105]<<11))-(0+(in_buffer[106]<<4)+(in_buffer[106]<<5)+(in_buffer[106]<<8)+(in_buffer[106]<<10))-(0+(in_buffer[107]<<1)+(in_buffer[107]<<3)+(in_buffer[107]<<7)+(in_buffer[107]<<10))+(0+(in_buffer[108]<<3)+(in_buffer[108]<<4)+(in_buffer[108]<<7)+(in_buffer[108]<<9))+(0-(in_buffer[109]<<1)-(in_buffer[109]<<4)+(in_buffer[109]<<7)+(in_buffer[109]<<11))+(0+(in_buffer[110]<<5)-(in_buffer[110]<<8)+(in_buffer[110]<<13))+(0+(in_buffer[111]<<1)+(in_buffer[111]<<2)-(in_buffer[111]<<8)+(in_buffer[111]<<10)+(in_buffer[111]<<11))-(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)-(in_buffer[112]<<5)+(in_buffer[112]<<8)-(in_buffer[112]<<10)+(in_buffer[112]<<13))-(0-(in_buffer[113]<<2)+(in_buffer[113]<<5)+(in_buffer[113]<<6)+(in_buffer[113]<<9)-(in_buffer[113]<<11)+(in_buffer[113]<<14))+(0+(in_buffer[114]<<0)+(in_buffer[114]<<2)-(in_buffer[114]<<4)-(in_buffer[114]<<7)+(in_buffer[114]<<11))+(0+(in_buffer[115]<<5)-(in_buffer[115]<<8)+(in_buffer[115]<<13))+(0-(in_buffer[116]<<1)+(in_buffer[116]<<4)-(in_buffer[116]<<6)+(in_buffer[116]<<8)+(in_buffer[116]<<9)+(in_buffer[116]<<12))-(0-(in_buffer[117]<<0)+(in_buffer[117]<<4)+(in_buffer[117]<<5)+(in_buffer[117]<<8)+(in_buffer[117]<<12))-(0-(in_buffer[118]<<0)+(in_buffer[118]<<3)-(in_buffer[118]<<6)+(in_buffer[118]<<10)+(in_buffer[118]<<12))+(0+(in_buffer[119]<<6)+(in_buffer[119]<<7)+(in_buffer[119]<<10)+(in_buffer[119]<<12))+(0-(in_buffer[120]<<0)-(in_buffer[120]<<3)+(in_buffer[120]<<8)+(in_buffer[120]<<11)+(in_buffer[120]<<12));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<3)-(in_buffer[0]<<5)+(in_buffer[0]<<8)+(in_buffer[0]<<9)+(in_buffer[0]<<12)+(in_buffer[0]<<13))-(0+(in_buffer[1]<<4)+(in_buffer[1]<<5)-(in_buffer[1]<<11)+(in_buffer[1]<<13)+(in_buffer[1]<<14))-(0-(in_buffer[2]<<2)+(in_buffer[2]<<4)+(in_buffer[2]<<5)+(in_buffer[2]<<11)+(in_buffer[2]<<15))-(0+(in_buffer[3]<<2)-(in_buffer[3]<<4)-(in_buffer[3]<<7)+(in_buffer[3]<<10)+(in_buffer[3]<<12))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<3)+(in_buffer[4]<<7)+(in_buffer[4]<<12))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<5)+(in_buffer[5]<<7)+(in_buffer[5]<<8))+(0-(in_buffer[6]<<1)+(in_buffer[6]<<11)+(in_buffer[6]<<12))+(0-(in_buffer[7]<<2)+(in_buffer[7]<<7)+(in_buffer[7]<<9)+(in_buffer[7]<<10))-(0-(in_buffer[8]<<0)-(in_buffer[8]<<3)+(in_buffer[8]<<6)+(in_buffer[8]<<9)+(in_buffer[8]<<11)+(in_buffer[8]<<13)+(in_buffer[8]<<15))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<5)+(in_buffer[9]<<8)+(in_buffer[9]<<11)+(in_buffer[9]<<15))-(0+(in_buffer[10]<<3)+(in_buffer[10]<<5)+(in_buffer[10]<<6)+(in_buffer[10]<<12)+(in_buffer[10]<<14))-(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)-(in_buffer[11]<<4)+(in_buffer[11]<<7)-(in_buffer[11]<<10)+(in_buffer[11]<<12)+(in_buffer[11]<<13))-(0-(in_buffer[12]<<4)-(in_buffer[12]<<7)+(in_buffer[12]<<10)+(in_buffer[12]<<14))-(0+(in_buffer[13]<<1)-(in_buffer[13]<<5)-(in_buffer[13]<<7)+(in_buffer[13]<<9)+(in_buffer[13]<<10)+(in_buffer[13]<<14))-(0-(in_buffer[14]<<1)-(in_buffer[14]<<4)+(in_buffer[14]<<9)+(in_buffer[14]<<12)+(in_buffer[14]<<13))+(0+(in_buffer[15]<<1)+(in_buffer[15]<<7)+(in_buffer[15]<<8)+(in_buffer[15]<<12))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<1)-(in_buffer[16]<<5)+(in_buffer[16]<<12))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<3)+(in_buffer[17]<<6)+(in_buffer[17]<<8)+(in_buffer[17]<<10)+(in_buffer[17]<<11))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)-(in_buffer[18]<<5)+(in_buffer[18]<<7)+(in_buffer[18]<<8)+(in_buffer[18]<<13))-(0+(in_buffer[19]<<2)-(in_buffer[19]<<6)-(in_buffer[19]<<11)+(in_buffer[19]<<14))-(0+(in_buffer[20]<<4)+(in_buffer[20]<<7)+(in_buffer[20]<<9)+(in_buffer[20]<<13)+(in_buffer[20]<<14))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<1)+(in_buffer[21]<<9)+(in_buffer[21]<<15))-(0-(in_buffer[22]<<0)+(in_buffer[22]<<4)-(in_buffer[22]<<7)-(in_buffer[22]<<10)+(in_buffer[22]<<13))-(0+(in_buffer[23]<<1)+(in_buffer[23]<<2)-(in_buffer[23]<<8)+(in_buffer[23]<<10)+(in_buffer[23]<<11))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)+(in_buffer[24]<<3)+(in_buffer[24]<<9)+(in_buffer[24]<<11))+(0+(in_buffer[25]<<1)-(in_buffer[25]<<4)+(in_buffer[25]<<9))+(0+(in_buffer[26]<<1)+(in_buffer[26]<<5)-(in_buffer[26]<<8)+(in_buffer[26]<<11))+(0+(in_buffer[27]<<0)+(in_buffer[27]<<4)-(in_buffer[27]<<7)+(in_buffer[27]<<10))+(0+(in_buffer[28]<<0)+(in_buffer[28]<<1)-(in_buffer[28]<<7)+(in_buffer[28]<<9)+(in_buffer[28]<<10))-(0+(in_buffer[29]<<3)+(in_buffer[29]<<4)+(in_buffer[29]<<7)+(in_buffer[29]<<9))+(0+(in_buffer[30]<<0)+(in_buffer[30]<<2)-(in_buffer[30]<<8)+(in_buffer[30]<<11)+(in_buffer[30]<<12))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<1)-(in_buffer[31]<<5)+(in_buffer[31]<<12))-(0+(in_buffer[32]<<0)+(in_buffer[32]<<2)+(in_buffer[32]<<4)+(in_buffer[32]<<6)-(in_buffer[32]<<9)+(in_buffer[32]<<12)+(in_buffer[32]<<15))-(0-(in_buffer[33]<<0)+(in_buffer[33]<<3)-(in_buffer[33]<<6)+(in_buffer[33]<<10)+(in_buffer[33]<<12))-(0-(in_buffer[34]<<0)+(in_buffer[34]<<3)-(in_buffer[34]<<5)+(in_buffer[34]<<7)+(in_buffer[34]<<8)+(in_buffer[34]<<11))+(0+(in_buffer[35]<<0)+(in_buffer[35]<<2)+(in_buffer[35]<<5)+(in_buffer[35]<<7)+(in_buffer[35]<<10)+(in_buffer[35]<<11))-(0-(in_buffer[36]<<0)+(in_buffer[36]<<5)+(in_buffer[36]<<6)-(in_buffer[36]<<9)+(in_buffer[36]<<11)+(in_buffer[36]<<12))-(0-(in_buffer[37]<<1)+(in_buffer[37]<<6)+(in_buffer[37]<<8)+(in_buffer[37]<<9))-(0+(in_buffer[38]<<0)+(in_buffer[38]<<3)-(in_buffer[38]<<5)-(in_buffer[38]<<8)-(in_buffer[38]<<10)+(in_buffer[38]<<13))-(0-(in_buffer[39]<<0)+(in_buffer[39]<<2)+(in_buffer[39]<<3)+(in_buffer[39]<<6)+(in_buffer[39]<<8)+(in_buffer[39]<<10)+(in_buffer[39]<<11))-(0+(in_buffer[40]<<2)+(in_buffer[40]<<4)+(in_buffer[40]<<8)+(in_buffer[40]<<11))+(0+(in_buffer[41]<<5)+(in_buffer[41]<<6)+(in_buffer[41]<<9)+(in_buffer[41]<<11))+(0+(in_buffer[42]<<0)+(in_buffer[42]<<6)+(in_buffer[42]<<7)+(in_buffer[42]<<11))-(0+(in_buffer[43]<<1)+(in_buffer[43]<<3)-(in_buffer[43]<<5)-(in_buffer[43]<<8)+(in_buffer[43]<<12))-(0-(in_buffer[44]<<1)+(in_buffer[44]<<6)+(in_buffer[44]<<8)+(in_buffer[44]<<9))+(0-(in_buffer[45]<<0)-(in_buffer[45]<<2)-(in_buffer[45]<<4)+(in_buffer[45]<<8)+(in_buffer[45]<<9))+(0-(in_buffer[46]<<1)+(in_buffer[46]<<5)-(in_buffer[46]<<7)-(in_buffer[46]<<9)+(in_buffer[46]<<12))-(0+(in_buffer[47]<<0)+(in_buffer[47]<<1)-(in_buffer[47]<<7)+(in_buffer[47]<<9)+(in_buffer[47]<<10))-(0-(in_buffer[48]<<0)+(in_buffer[48]<<5)+(in_buffer[48]<<7)+(in_buffer[48]<<8))-(0+(in_buffer[49]<<2)-(in_buffer[49]<<4)-(in_buffer[49]<<7)+(in_buffer[49]<<10)+(in_buffer[49]<<12))-(0-(in_buffer[50]<<0)+(in_buffer[50]<<3)+(in_buffer[50]<<4)+(in_buffer[50]<<7)-(in_buffer[50]<<9)+(in_buffer[50]<<12))-(0+(in_buffer[51]<<0)+(in_buffer[51]<<1)+(in_buffer[51]<<4)+(in_buffer[51]<<6))+(0+(in_buffer[52]<<0)+(in_buffer[52]<<6)+(in_buffer[52]<<7)+(in_buffer[52]<<11))+(0-(in_buffer[53]<<0)+(in_buffer[53]<<3)-(in_buffer[53]<<5)+(in_buffer[53]<<7)+(in_buffer[53]<<8)+(in_buffer[53]<<11))+(0+(in_buffer[54]<<0)-(in_buffer[54]<<2)-(in_buffer[54]<<5)+(in_buffer[54]<<8)+(in_buffer[54]<<10))-(0-(in_buffer[55]<<0)+(in_buffer[55]<<4)-(in_buffer[55]<<7)-(in_buffer[55]<<10)+(in_buffer[55]<<13))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<1)+(in_buffer[56]<<4)+(in_buffer[56]<<6))+(0+(in_buffer[57]<<0)+(in_buffer[57]<<3)+(in_buffer[57]<<5)+(in_buffer[57]<<9)+(in_buffer[57]<<10))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<1)+(in_buffer[58]<<4)+(in_buffer[58]<<6))+(0-(in_buffer[59]<<1)+(in_buffer[59]<<6)+(in_buffer[59]<<8)+(in_buffer[59]<<9))-(0+(in_buffer[60]<<2)+(in_buffer[60]<<3)+(in_buffer[60]<<6)+(in_buffer[60]<<8))-(0+(in_buffer[61]<<0)-(in_buffer[61]<<3)+(in_buffer[61]<<8))+(0+(in_buffer[62]<<1)+(in_buffer[62]<<3)+(in_buffer[62]<<7)+(in_buffer[62]<<10))+(0+(in_buffer[63]<<0)+(in_buffer[63]<<1)-(in_buffer[63]<<7)+(in_buffer[63]<<9)+(in_buffer[63]<<10))-(0+(in_buffer[64]<<0)+(in_buffer[64]<<1)-(in_buffer[64]<<7)+(in_buffer[64]<<9)+(in_buffer[64]<<10))+(0+(in_buffer[65]<<1)+(in_buffer[65]<<5)-(in_buffer[65]<<8)+(in_buffer[65]<<11))-(0-(in_buffer[66]<<0)+(in_buffer[66]<<5)+(in_buffer[66]<<6)-(in_buffer[66]<<9)+(in_buffer[66]<<11)+(in_buffer[66]<<12))-(0+(in_buffer[67]<<5)-(in_buffer[67]<<8)+(in_buffer[67]<<13))+(0-(in_buffer[68]<<1)-(in_buffer[68]<<3)-(in_buffer[68]<<5)+(in_buffer[68]<<9)+(in_buffer[68]<<10))+(0-(in_buffer[69]<<0)+(in_buffer[69]<<2)+(in_buffer[69]<<3)+(in_buffer[69]<<6)+(in_buffer[69]<<8)+(in_buffer[69]<<10)+(in_buffer[69]<<11))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<2)+(in_buffer[70]<<3)+(in_buffer[70]<<9)+(in_buffer[70]<<11))+(0-(in_buffer[71]<<0)-(in_buffer[71]<<2)+(in_buffer[71]<<5)+(in_buffer[71]<<11))+(0+(in_buffer[72]<<1)+(in_buffer[72]<<2)+(in_buffer[72]<<5)+(in_buffer[72]<<7))+(0-(in_buffer[73]<<1)-(in_buffer[73]<<3)-(in_buffer[73]<<5)+(in_buffer[73]<<9)+(in_buffer[73]<<10))-(0+(in_buffer[75]<<4)+(in_buffer[75]<<5)+(in_buffer[75]<<8)+(in_buffer[75]<<10))+(0+(in_buffer[76]<<0)+(in_buffer[76]<<1)-(in_buffer[76]<<4)-(in_buffer[76]<<6)-(in_buffer[76]<<8)+(in_buffer[76]<<10)+(in_buffer[76]<<11))+(0-(in_buffer[77]<<0)-(in_buffer[77]<<3)+(in_buffer[77]<<6)+(in_buffer[77]<<10))-(0-(in_buffer[78]<<4)+(in_buffer[78]<<9)+(in_buffer[78]<<11)+(in_buffer[78]<<12))+(0+(in_buffer[79]<<3)-(in_buffer[79]<<6)+(in_buffer[79]<<11))+(0+(in_buffer[80]<<1)+(in_buffer[80]<<4)+(in_buffer[80]<<6)+(in_buffer[80]<<10)+(in_buffer[80]<<11))-(0+(in_buffer[81]<<2)+(in_buffer[81]<<3)+(in_buffer[81]<<6)+(in_buffer[81]<<8))+(0-(in_buffer[82]<<1)-(in_buffer[82]<<3)-(in_buffer[82]<<5)+(in_buffer[82]<<9)+(in_buffer[82]<<10))-(0+(in_buffer[83]<<0)+(in_buffer[83]<<1)+(in_buffer[83]<<4)+(in_buffer[83]<<6))+(0+(in_buffer[84]<<0)-(in_buffer[84]<<2)-(in_buffer[84]<<5)+(in_buffer[84]<<8)+(in_buffer[84]<<10))+(0+(in_buffer[85]<<0)-(in_buffer[85]<<3)+(in_buffer[85]<<8))+(0+(in_buffer[86]<<1)+(in_buffer[86]<<2)+(in_buffer[86]<<5)+(in_buffer[86]<<7))+(0+(in_buffer[87]<<0)-(in_buffer[87]<<2)+(in_buffer[87]<<5)+(in_buffer[87]<<7)+(in_buffer[87]<<8)+(in_buffer[87]<<11)+(in_buffer[87]<<12))+(0+(in_buffer[88]<<1)+(in_buffer[88]<<2)-(in_buffer[88]<<8)+(in_buffer[88]<<10)+(in_buffer[88]<<11))+(0-(in_buffer[89]<<0)+(in_buffer[89]<<3)+(in_buffer[89]<<4)+(in_buffer[89]<<7)-(in_buffer[89]<<9)+(in_buffer[89]<<12))+(0+(in_buffer[90]<<0)+(in_buffer[90]<<2)-(in_buffer[90]<<4)-(in_buffer[90]<<7)+(in_buffer[90]<<11))-(0+(in_buffer[91]<<2)+(in_buffer[91]<<3)+(in_buffer[91]<<6)+(in_buffer[91]<<8))-(0-(in_buffer[92]<<0)+(in_buffer[92]<<4)-(in_buffer[92]<<6)-(in_buffer[92]<<8)+(in_buffer[92]<<11))+(0+(in_buffer[93]<<0)+(in_buffer[93]<<3)+(in_buffer[93]<<5)+(in_buffer[93]<<9)+(in_buffer[93]<<10))+(0-(in_buffer[94]<<2)+(in_buffer[94]<<7)+(in_buffer[94]<<9)+(in_buffer[94]<<10))+(0+(in_buffer[95]<<3)+(in_buffer[95]<<4)+(in_buffer[95]<<7)+(in_buffer[95]<<9))-(0+(in_buffer[96]<<0)+(in_buffer[96]<<6)+(in_buffer[96]<<7)+(in_buffer[96]<<11))+(0+(in_buffer[97]<<2)-(in_buffer[97]<<5)+(in_buffer[97]<<10))+(0-(in_buffer[98]<<1)+(in_buffer[98]<<5)-(in_buffer[98]<<7)-(in_buffer[98]<<9)+(in_buffer[98]<<12))-(0-(in_buffer[99]<<1)+(in_buffer[99]<<4)-(in_buffer[99]<<6)+(in_buffer[99]<<8)+(in_buffer[99]<<9)+(in_buffer[99]<<12))+(0+(in_buffer[100]<<0)+(in_buffer[100]<<2)-(in_buffer[100]<<8)+(in_buffer[100]<<11)+(in_buffer[100]<<12))-(0-(in_buffer[101]<<2)-(in_buffer[101]<<4)-(in_buffer[101]<<6)+(in_buffer[101]<<10)+(in_buffer[101]<<11))-(0+(in_buffer[102]<<1)+(in_buffer[102]<<3)-(in_buffer[102]<<5)-(in_buffer[102]<<8)+(in_buffer[102]<<12))+(0+(in_buffer[103]<<0)+(in_buffer[103]<<1)-(in_buffer[103]<<5)+(in_buffer[103]<<12))+(0+(in_buffer[104]<<2)-(in_buffer[104]<<4)-(in_buffer[104]<<7)+(in_buffer[104]<<10)+(in_buffer[104]<<12))+(0-(in_buffer[105]<<2)+(in_buffer[105]<<6)-(in_buffer[105]<<8)-(in_buffer[105]<<10)+(in_buffer[105]<<13))-(0+(in_buffer[106]<<0)+(in_buffer[106]<<1)+(in_buffer[106]<<4)+(in_buffer[106]<<6))-(0+(in_buffer[107]<<2)+(in_buffer[107]<<4)+(in_buffer[107]<<8)+(in_buffer[107]<<11))+(0+(in_buffer[108]<<0)+(in_buffer[108]<<3)+(in_buffer[108]<<5)+(in_buffer[108]<<9)+(in_buffer[108]<<10))+(0+(in_buffer[109]<<2)+(in_buffer[109]<<4)+(in_buffer[109]<<8)+(in_buffer[109]<<11))+(0-(in_buffer[110]<<0)+(in_buffer[110]<<3)+(in_buffer[110]<<5)-(in_buffer[110]<<9)+(in_buffer[110]<<13))+(0+(in_buffer[111]<<0)+(in_buffer[111]<<1)-(in_buffer[111]<<7)+(in_buffer[111]<<9)+(in_buffer[111]<<10))-(0-(in_buffer[112]<<0)+(in_buffer[112]<<10)+(in_buffer[112]<<11))+(0-(in_buffer[113]<<4)+(in_buffer[113]<<9)+(in_buffer[113]<<11)+(in_buffer[113]<<12))+(0+(in_buffer[114]<<1)+(in_buffer[114]<<3)+(in_buffer[114]<<7)+(in_buffer[114]<<10))-(0+(in_buffer[115]<<0)+(in_buffer[115]<<2)-(in_buffer[115]<<4)-(in_buffer[115]<<7)+(in_buffer[115]<<11))+(0+(in_buffer[116]<<0)+(in_buffer[116]<<1)+(in_buffer[116]<<4)+(in_buffer[116]<<6))+(0-(in_buffer[117]<<0)+(in_buffer[117]<<4)+(in_buffer[117]<<5)+(in_buffer[117]<<8)+(in_buffer[117]<<12))+(0+(in_buffer[118]<<0)+(in_buffer[118]<<4)-(in_buffer[118]<<7)+(in_buffer[118]<<10))+(0+(in_buffer[119]<<0)+(in_buffer[119]<<2)-(in_buffer[119]<<4)-(in_buffer[119]<<7)+(in_buffer[119]<<11))+(0-(in_buffer[120]<<1)+(in_buffer[120]<<4)-(in_buffer[120]<<7)+(in_buffer[120]<<11)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0-(0+(in_buffer[0]<<1)+(in_buffer[0]<<3)+(in_buffer[0]<<6)+(in_buffer[0]<<8)+(in_buffer[0]<<11)+(in_buffer[0]<<12))-(0-(in_buffer[1]<<2)-(in_buffer[1]<<5)+(in_buffer[1]<<8)+(in_buffer[1]<<12))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<2)+(in_buffer[2]<<5)+(in_buffer[2]<<7))-(0-(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<4)+(in_buffer[3]<<7)-(in_buffer[3]<<9)+(in_buffer[3]<<12))-(0+(in_buffer[4]<<0)-(in_buffer[4]<<4)-(in_buffer[4]<<9)+(in_buffer[4]<<12))+(0-(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<5)+(in_buffer[5]<<11))-(0-(in_buffer[6]<<0)-(in_buffer[6]<<3)+(in_buffer[6]<<8)+(in_buffer[6]<<11)+(in_buffer[6]<<12))-(0+(in_buffer[7]<<0)-(in_buffer[7]<<2)-(in_buffer[7]<<4)+(in_buffer[7]<<7)+(in_buffer[7]<<10)+(in_buffer[7]<<12))-(0-(in_buffer[8]<<1)+(in_buffer[8]<<3)+(in_buffer[8]<<4)+(in_buffer[8]<<7)+(in_buffer[8]<<9)+(in_buffer[8]<<11)+(in_buffer[8]<<12))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<6)+(in_buffer[9]<<9))+(0+(in_buffer[10]<<2)+(in_buffer[10]<<3)+(in_buffer[10]<<6)+(in_buffer[10]<<8))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3)-(in_buffer[11]<<6)-(in_buffer[11]<<8)+(in_buffer[11]<<13))-(0+(in_buffer[12]<<1)-(in_buffer[12]<<5)-(in_buffer[12]<<10)+(in_buffer[12]<<13))-(0-(in_buffer[13]<<1)-(in_buffer[13]<<3)+(in_buffer[13]<<6)+(in_buffer[13]<<12))+(0-(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<5)+(in_buffer[14]<<11))-(0-(in_buffer[15]<<0)-(in_buffer[15]<<3)+(in_buffer[15]<<6)+(in_buffer[15]<<10))-(0-(in_buffer[16]<<1)-(in_buffer[16]<<3)-(in_buffer[16]<<5)+(in_buffer[16]<<9)+(in_buffer[16]<<10))+(0+(in_buffer[17]<<2)-(in_buffer[17]<<5)+(in_buffer[17]<<10))+(0-(in_buffer[18]<<0)+(in_buffer[18]<<4)+(in_buffer[18]<<5)+(in_buffer[18]<<8)+(in_buffer[18]<<12))-(0-(in_buffer[19]<<1)-(in_buffer[19]<<3)-(in_buffer[19]<<5)+(in_buffer[19]<<9)+(in_buffer[19]<<10))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<3)+(in_buffer[20]<<7)+(in_buffer[20]<<9)+(in_buffer[20]<<11)+(in_buffer[20]<<13))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)-(in_buffer[21]<<6)-(in_buffer[21]<<10)+(in_buffer[21]<<12)+(in_buffer[21]<<13))-(0+(in_buffer[22]<<2)+(in_buffer[22]<<6)-(in_buffer[22]<<9)+(in_buffer[22]<<12))-(0-(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<7)+(in_buffer[23]<<9)+(in_buffer[23]<<12))-(0-(in_buffer[24]<<1)-(in_buffer[24]<<3)-(in_buffer[24]<<5)+(in_buffer[24]<<9)+(in_buffer[24]<<10))-(0+(in_buffer[25]<<2)+(in_buffer[25]<<3)+(in_buffer[25]<<6)+(in_buffer[25]<<8))+(0+(in_buffer[26]<<0)+(in_buffer[26]<<1)+(in_buffer[26]<<4)+(in_buffer[26]<<6))-(0+(in_buffer[27]<<0)+(in_buffer[27]<<6)+(in_buffer[27]<<7)+(in_buffer[27]<<11))-(0+(in_buffer[28]<<3)+(in_buffer[28]<<4)+(in_buffer[28]<<7)+(in_buffer[28]<<9))+(0-(in_buffer[29]<<0)+(in_buffer[29]<<4)-(in_buffer[29]<<6)-(in_buffer[29]<<8)+(in_buffer[29]<<11))+(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)-(in_buffer[30]<<4)+(in_buffer[30]<<8)+(in_buffer[30]<<9))-(0-(in_buffer[31]<<1)+(in_buffer[31]<<5)-(in_buffer[31]<<7)-(in_buffer[31]<<9)+(in_buffer[31]<<12))+(0-(in_buffer[32]<<1)-(in_buffer[32]<<3)+(in_buffer[32]<<6)+(in_buffer[32]<<12))+(0+(in_buffer[33]<<3)+(in_buffer[33]<<4)+(in_buffer[33]<<7)+(in_buffer[33]<<9))-(0+(in_buffer[34]<<4)+(in_buffer[34]<<5)+(in_buffer[34]<<8)+(in_buffer[34]<<10))-(0+(in_buffer[35]<<2)-(in_buffer[35]<<5)+(in_buffer[35]<<10))-(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)-(in_buffer[36]<<4)+(in_buffer[36]<<8)+(in_buffer[36]<<9))-(0+(in_buffer[37]<<4)+(in_buffer[37]<<5)+(in_buffer[37]<<8)+(in_buffer[37]<<10))-(0+(in_buffer[38]<<0)+(in_buffer[38]<<3)+(in_buffer[38]<<7)+(in_buffer[38]<<12))-(0+(in_buffer[40]<<3)+(in_buffer[40]<<4)+(in_buffer[40]<<7)+(in_buffer[40]<<9))-(0-(in_buffer[41]<<1)-(in_buffer[41]<<3)-(in_buffer[41]<<5)+(in_buffer[41]<<9)+(in_buffer[41]<<10))+(0+(in_buffer[42]<<4)-(in_buffer[42]<<7)+(in_buffer[42]<<12))+(0-(in_buffer[43]<<1)+(in_buffer[43]<<11)+(in_buffer[43]<<12))+(0+(in_buffer[44]<<1)+(in_buffer[44]<<4)+(in_buffer[44]<<6)+(in_buffer[44]<<10)+(in_buffer[44]<<11))+(0-(in_buffer[45]<<0)+(in_buffer[45]<<3)-(in_buffer[45]<<5)+(in_buffer[45]<<7)+(in_buffer[45]<<8)+(in_buffer[45]<<11))+(0+(in_buffer[46]<<0)+(in_buffer[46]<<2)+(in_buffer[46]<<5)+(in_buffer[46]<<7)+(in_buffer[46]<<10)+(in_buffer[46]<<11))+(0+(in_buffer[47]<<4)-(in_buffer[47]<<7)+(in_buffer[47]<<12))+(0+(in_buffer[48]<<4)+(in_buffer[48]<<5)+(in_buffer[48]<<8)+(in_buffer[48]<<10))+(0-(in_buffer[49]<<0)+(in_buffer[49]<<3)-(in_buffer[49]<<5)+(in_buffer[49]<<7)+(in_buffer[49]<<8)+(in_buffer[49]<<11))+(0+(in_buffer[50]<<0)+(in_buffer[50]<<2)+(in_buffer[50]<<6)+(in_buffer[50]<<9))+(0-(in_buffer[51]<<0)+(in_buffer[51]<<4)-(in_buffer[51]<<6)-(in_buffer[51]<<8)+(in_buffer[51]<<11))+(0+(in_buffer[52]<<3)+(in_buffer[52]<<4)+(in_buffer[52]<<7)+(in_buffer[52]<<9))+(0+(in_buffer[54]<<1)+(in_buffer[54]<<3)+(in_buffer[54]<<6)+(in_buffer[54]<<8)+(in_buffer[54]<<11)+(in_buffer[54]<<12))-(0+(in_buffer[55]<<1)+(in_buffer[55]<<3)-(in_buffer[55]<<5)-(in_buffer[55]<<8)+(in_buffer[55]<<12))-(0+(in_buffer[56]<<2)-(in_buffer[56]<<5)+(in_buffer[56]<<10))+(0-(in_buffer[57]<<0)+(in_buffer[57]<<4)-(in_buffer[57]<<6)-(in_buffer[57]<<8)+(in_buffer[57]<<11))+(0+(in_buffer[58]<<2)+(in_buffer[58]<<5)+(in_buffer[58]<<7)+(in_buffer[58]<<11)+(in_buffer[58]<<12))+(0-(in_buffer[60]<<0)+(in_buffer[60]<<3)+(in_buffer[60]<<4)+(in_buffer[60]<<7)-(in_buffer[60]<<9)+(in_buffer[60]<<12))+(0+(in_buffer[61]<<3)+(in_buffer[61]<<4)+(in_buffer[61]<<7)+(in_buffer[61]<<9))+(0-(in_buffer[62]<<0)+(in_buffer[62]<<3)-(in_buffer[62]<<6)+(in_buffer[62]<<10)+(in_buffer[62]<<12))+(0-(in_buffer[63]<<2)-(in_buffer[63]<<4)-(in_buffer[63]<<6)+(in_buffer[63]<<10)+(in_buffer[63]<<11))+(0-(in_buffer[64]<<0)+(in_buffer[64]<<3)+(in_buffer[64]<<4)+(in_buffer[64]<<7)-(in_buffer[64]<<9)+(in_buffer[64]<<12))+(0+(in_buffer[65]<<2)-(in_buffer[65]<<4)-(in_buffer[65]<<7)+(in_buffer[65]<<10)+(in_buffer[65]<<12))+(0+(in_buffer[66]<<1)+(in_buffer[66]<<4)+(in_buffer[66]<<6)+(in_buffer[66]<<10)+(in_buffer[66]<<11))-(0-(in_buffer[67]<<1)-(in_buffer[67]<<4)+(in_buffer[67]<<7)+(in_buffer[67]<<11))-(0-(in_buffer[68]<<0)+(in_buffer[68]<<4)-(in_buffer[68]<<6)-(in_buffer[68]<<8)+(in_buffer[68]<<11))+(0+(in_buffer[69]<<6)+(in_buffer[69]<<7)+(in_buffer[69]<<10)+(in_buffer[69]<<12))+(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)-(in_buffer[70]<<4)+(in_buffer[70]<<8)+(in_buffer[70]<<9))+(0+(in_buffer[71]<<0)+(in_buffer[71]<<6)+(in_buffer[71]<<7)+(in_buffer[71]<<11))+(0+(in_buffer[72]<<0)+(in_buffer[72]<<2)+(in_buffer[72]<<6)+(in_buffer[72]<<9))+(0+(in_buffer[73]<<0)-(in_buffer[73]<<2)-(in_buffer[73]<<4)+(in_buffer[73]<<7)+(in_buffer[73]<<10)+(in_buffer[73]<<12))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<2)-(in_buffer[74]<<5)+(in_buffer[74]<<8)+(in_buffer[74]<<10))+(0+(in_buffer[75]<<0)+(in_buffer[75]<<2)-(in_buffer[75]<<4)-(in_buffer[75]<<7)+(in_buffer[75]<<11))-(0+(in_buffer[76]<<0)+(in_buffer[76]<<1)+(in_buffer[76]<<4)+(in_buffer[76]<<6))+(0+(in_buffer[77]<<0)+(in_buffer[77]<<1)+(in_buffer[77]<<4)+(in_buffer[77]<<8)+(in_buffer[77]<<10)+(in_buffer[77]<<12))-(0+(in_buffer[78]<<2)+(in_buffer[78]<<6)-(in_buffer[78]<<9)+(in_buffer[78]<<12))-(0+(in_buffer[79]<<0)+(in_buffer[79]<<1)-(in_buffer[79]<<5)+(in_buffer[79]<<12))+(0+(in_buffer[80]<<2)+(in_buffer[80]<<3)+(in_buffer[80]<<6)+(in_buffer[80]<<8))-(0+(in_buffer[81]<<0)+(in_buffer[81]<<6)+(in_buffer[81]<<7)+(in_buffer[81]<<11))+(0+(in_buffer[82]<<2)-(in_buffer[82]<<4)-(in_buffer[82]<<7)+(in_buffer[82]<<10)+(in_buffer[82]<<12))+(0-(in_buffer[83]<<0)-(in_buffer[83]<<2)+(in_buffer[83]<<5)+(in_buffer[83]<<11))+(0-(in_buffer[84]<<1)-(in_buffer[84]<<3)+(in_buffer[84]<<6)+(in_buffer[84]<<12))-(0+(in_buffer[85]<<0)+(in_buffer[85]<<1)+(in_buffer[85]<<4)+(in_buffer[85]<<6))-(0+(in_buffer[86]<<1)+(in_buffer[86]<<7)+(in_buffer[86]<<8)+(in_buffer[86]<<12))+(0+(in_buffer[87]<<0)-(in_buffer[87]<<3)-(in_buffer[87]<<5)-(in_buffer[87]<<7)+(in_buffer[87]<<10)+(in_buffer[87]<<11))+(0-(in_buffer[88]<<2)+(in_buffer[88]<<7)+(in_buffer[88]<<9)+(in_buffer[88]<<10))+(0+(in_buffer[89]<<0)-(in_buffer[89]<<3)+(in_buffer[89]<<8))-(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)-(in_buffer[90]<<4)+(in_buffer[90]<<8)+(in_buffer[90]<<9))-(0-(in_buffer[91]<<1)+(in_buffer[91]<<6)+(in_buffer[91]<<8)+(in_buffer[91]<<9))-(0+(in_buffer[92]<<0)+(in_buffer[92]<<5)+(in_buffer[92]<<8)+(in_buffer[92]<<9)+(in_buffer[92]<<12))+(0-(in_buffer[93]<<1)-(in_buffer[93]<<3)+(in_buffer[93]<<6)+(in_buffer[93]<<12))+(0-(in_buffer[94]<<0)-(in_buffer[94]<<2)+(in_buffer[94]<<7)+(in_buffer[94]<<9)+(in_buffer[94]<<12))+(0+(in_buffer[95]<<0)+(in_buffer[95]<<1)-(in_buffer[95]<<4)-(in_buffer[95]<<6)-(in_buffer[95]<<8)+(in_buffer[95]<<10)+(in_buffer[95]<<11))-(0+(in_buffer[96]<<0)+(in_buffer[96]<<4)-(in_buffer[96]<<7)+(in_buffer[96]<<10))-(0-(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<7)+(in_buffer[97]<<9)+(in_buffer[97]<<12))+(0+(in_buffer[98]<<2)+(in_buffer[98]<<3)+(in_buffer[98]<<6)+(in_buffer[98]<<8))-(0+(in_buffer[99]<<0)+(in_buffer[99]<<3)+(in_buffer[99]<<5)+(in_buffer[99]<<9)+(in_buffer[99]<<10))+(0-(in_buffer[100]<<0)-(in_buffer[100]<<2)-(in_buffer[100]<<5)+(in_buffer[100]<<8)-(in_buffer[100]<<10)+(in_buffer[100]<<13))+(0+(in_buffer[101]<<0)+(in_buffer[101]<<4)+(in_buffer[101]<<6)+(in_buffer[101]<<11)+(in_buffer[101]<<12))+(0-(in_buffer[102]<<0)+(in_buffer[102]<<4)-(in_buffer[102]<<6)-(in_buffer[102]<<8)+(in_buffer[102]<<11))-(0-(in_buffer[103]<<0)+(in_buffer[103]<<10)+(in_buffer[103]<<11))+(0+(in_buffer[104]<<4)+(in_buffer[104]<<5)+(in_buffer[104]<<8)+(in_buffer[104]<<10))+(0+(in_buffer[105]<<0)-(in_buffer[105]<<2)-(in_buffer[105]<<5)+(in_buffer[105]<<8)+(in_buffer[105]<<10))+(0+(in_buffer[106]<<4)-(in_buffer[106]<<7)+(in_buffer[106]<<12))+(0+(in_buffer[107]<<3)+(in_buffer[107]<<5)+(in_buffer[107]<<9)+(in_buffer[107]<<12))+(0+(in_buffer[108]<<0)+(in_buffer[108]<<1)-(in_buffer[108]<<4)-(in_buffer[108]<<6)-(in_buffer[108]<<8)+(in_buffer[108]<<10)+(in_buffer[108]<<11))-(0-(in_buffer[109]<<3)-(in_buffer[109]<<5)-(in_buffer[109]<<7)+(in_buffer[109]<<11)+(in_buffer[109]<<12))+(0-(in_buffer[110]<<0)-(in_buffer[110]<<2)+(in_buffer[110]<<5)+(in_buffer[110]<<11))+(0+(in_buffer[111]<<0)+(in_buffer[111]<<2)+(in_buffer[111]<<3)-(in_buffer[111]<<6)-(in_buffer[111]<<8)+(in_buffer[111]<<13))+(0+(in_buffer[112]<<2)+(in_buffer[112]<<3)+(in_buffer[112]<<6)+(in_buffer[112]<<8))-(0-(in_buffer[113]<<3)+(in_buffer[113]<<8)+(in_buffer[113]<<10)+(in_buffer[113]<<11))-(0-(in_buffer[114]<<2)+(in_buffer[114]<<7)+(in_buffer[114]<<9)+(in_buffer[114]<<10))+(0-(in_buffer[115]<<0)+(in_buffer[115]<<4)-(in_buffer[115]<<6)-(in_buffer[115]<<8)+(in_buffer[115]<<11))-(0-(in_buffer[116]<<0)+(in_buffer[116]<<10)+(in_buffer[116]<<11))-(0+(in_buffer[117]<<5)+(in_buffer[117]<<6)+(in_buffer[117]<<9)+(in_buffer[117]<<11))-(0+(in_buffer[118]<<0)+(in_buffer[118]<<4)+(in_buffer[118]<<6)+(in_buffer[118]<<11)+(in_buffer[118]<<12))-(0+(in_buffer[119]<<1)+(in_buffer[119]<<3)+(in_buffer[119]<<7)+(in_buffer[119]<<10))-(0-(in_buffer[120]<<0)+(in_buffer[120]<<3)-(in_buffer[120]<<6)+(in_buffer[120]<<10)+(in_buffer[120]<<12));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight10;
assign in_buffer_weight10=0-(0+(in_buffer[0]<<3)+(in_buffer[0]<<4)+(in_buffer[0]<<7)+(in_buffer[0]<<9))-(0-(in_buffer[1]<<1)-(in_buffer[1]<<4)-(in_buffer[1]<<6)-(in_buffer[1]<<8)+(in_buffer[1]<<11)+(in_buffer[1]<<14))-(0+(in_buffer[2]<<2)+(in_buffer[2]<<8)+(in_buffer[2]<<9)+(in_buffer[2]<<13))-(0+(in_buffer[3]<<3)-(in_buffer[3]<<6)+(in_buffer[3]<<11))+(0-(in_buffer[4]<<0)+(in_buffer[4]<<5)+(in_buffer[4]<<7)+(in_buffer[4]<<8))-(0-(in_buffer[5]<<1)+(in_buffer[5]<<5)-(in_buffer[5]<<7)-(in_buffer[5]<<9)+(in_buffer[5]<<12))+(0+(in_buffer[6]<<5)+(in_buffer[6]<<6)+(in_buffer[6]<<9)+(in_buffer[6]<<11))+(0-(in_buffer[7]<<2)+(in_buffer[7]<<7)+(in_buffer[7]<<9)+(in_buffer[7]<<10))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<4)+(in_buffer[8]<<8)+(in_buffer[8]<<11))-(0-(in_buffer[9]<<0)-(in_buffer[9]<<4)-(in_buffer[9]<<6)-(in_buffer[9]<<8)-(in_buffer[9]<<10)+(in_buffer[9]<<14))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<3)+(in_buffer[10]<<5)-(in_buffer[10]<<7)+(in_buffer[10]<<10)+(in_buffer[10]<<13))-(0-(in_buffer[11]<<3)+(in_buffer[11]<<7)-(in_buffer[11]<<9)-(in_buffer[11]<<11)+(in_buffer[11]<<14))+(0+(in_buffer[12]<<1)+(in_buffer[12]<<7)+(in_buffer[12]<<8)+(in_buffer[12]<<12))+(0+(in_buffer[13]<<0)-(in_buffer[13]<<2)-(in_buffer[13]<<5)+(in_buffer[13]<<8)+(in_buffer[13]<<10))-(0-(in_buffer[14]<<3)+(in_buffer[14]<<8)+(in_buffer[14]<<10)+(in_buffer[14]<<11))+(0-(in_buffer[15]<<1)-(in_buffer[15]<<4)+(in_buffer[15]<<7)+(in_buffer[15]<<11))-(0+(in_buffer[16]<<4)+(in_buffer[16]<<5)+(in_buffer[16]<<8)+(in_buffer[16]<<10))+(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)+(in_buffer[17]<<5)+(in_buffer[17]<<11))-(0+(in_buffer[18]<<0)-(in_buffer[18]<<3)+(in_buffer[18]<<8))+(0+(in_buffer[19]<<5)+(in_buffer[19]<<6)+(in_buffer[19]<<9)+(in_buffer[19]<<11))+(0+(in_buffer[20]<<2)-(in_buffer[20]<<4)+(in_buffer[20]<<8)-(in_buffer[20]<<10)+(in_buffer[20]<<14))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<5)+(in_buffer[21]<<8)-(in_buffer[21]<<11)+(in_buffer[21]<<13)+(in_buffer[21]<<14))-(0+(in_buffer[22]<<0)-(in_buffer[22]<<2)-(in_buffer[22]<<4)+(in_buffer[22]<<7)+(in_buffer[22]<<10)+(in_buffer[22]<<12))+(0-(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<4)+(in_buffer[23]<<7)+(in_buffer[23]<<9)+(in_buffer[23]<<11)+(in_buffer[23]<<12))+(0+(in_buffer[24]<<0)-(in_buffer[24]<<3)-(in_buffer[24]<<6)-(in_buffer[24]<<9)+(in_buffer[24]<<11)+(in_buffer[24]<<12))-(0+(in_buffer[25]<<1)+(in_buffer[25]<<5)-(in_buffer[25]<<8)+(in_buffer[25]<<11))-(0-(in_buffer[26]<<0)+(in_buffer[26]<<5)+(in_buffer[26]<<6)-(in_buffer[26]<<9)+(in_buffer[26]<<11)+(in_buffer[26]<<12))-(0+(in_buffer[27]<<0)+(in_buffer[27]<<2)+(in_buffer[27]<<4)-(in_buffer[27]<<6)+(in_buffer[27]<<9)+(in_buffer[27]<<12))+(0+(in_buffer[28]<<4)+(in_buffer[28]<<5)+(in_buffer[28]<<8)+(in_buffer[28]<<10))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<1)+(in_buffer[29]<<4)+(in_buffer[29]<<6))+(0+(in_buffer[30]<<2)+(in_buffer[30]<<3)-(in_buffer[30]<<9)+(in_buffer[30]<<11)+(in_buffer[30]<<12))+(0-(in_buffer[31]<<1)+(in_buffer[31]<<6)+(in_buffer[31]<<7)-(in_buffer[31]<<10)+(in_buffer[31]<<12)+(in_buffer[31]<<13))-(0-(in_buffer[32]<<0)+(in_buffer[32]<<5)+(in_buffer[32]<<6)-(in_buffer[32]<<9)+(in_buffer[32]<<11)+(in_buffer[32]<<12))-(0+(in_buffer[33]<<0)+(in_buffer[33]<<2)-(in_buffer[33]<<8)+(in_buffer[33]<<11)+(in_buffer[33]<<12))+(0-(in_buffer[34]<<1)+(in_buffer[34]<<6)+(in_buffer[34]<<8)+(in_buffer[34]<<9))+(0-(in_buffer[35]<<0)+(in_buffer[35]<<4)+(in_buffer[35]<<5)+(in_buffer[35]<<8)+(in_buffer[35]<<12))-(0-(in_buffer[36]<<2)-(in_buffer[36]<<4)-(in_buffer[36]<<6)+(in_buffer[36]<<10)+(in_buffer[36]<<11))-(0+(in_buffer[37]<<2)+(in_buffer[37]<<5)+(in_buffer[37]<<7)+(in_buffer[37]<<11)+(in_buffer[37]<<12))-(0+(in_buffer[38]<<4)-(in_buffer[38]<<7)+(in_buffer[38]<<12))-(0+(in_buffer[39]<<2)+(in_buffer[39]<<3)+(in_buffer[39]<<6)+(in_buffer[39]<<8))-(0+(in_buffer[40]<<4)+(in_buffer[40]<<5)+(in_buffer[40]<<8)+(in_buffer[40]<<10))+(0-(in_buffer[41]<<1)-(in_buffer[41]<<3)+(in_buffer[41]<<6)+(in_buffer[41]<<12))+(0+(in_buffer[42]<<0)+(in_buffer[42]<<2)+(in_buffer[42]<<5)+(in_buffer[42]<<7)+(in_buffer[42]<<10)+(in_buffer[42]<<11))+(0+(in_buffer[43]<<3)+(in_buffer[43]<<4)+(in_buffer[43]<<7)+(in_buffer[43]<<9))-(0+(in_buffer[44]<<0)+(in_buffer[44]<<1)+(in_buffer[44]<<5)+(in_buffer[44]<<7)+(in_buffer[44]<<10)+(in_buffer[44]<<13))-(0+(in_buffer[45]<<2)+(in_buffer[45]<<5)+(in_buffer[45]<<7)+(in_buffer[45]<<11)+(in_buffer[45]<<12))+(0+(in_buffer[46]<<0)+(in_buffer[46]<<3)+(in_buffer[46]<<5)+(in_buffer[46]<<9)+(in_buffer[46]<<10))-(0+(in_buffer[47]<<0)-(in_buffer[47]<<3)-(in_buffer[47]<<5)-(in_buffer[47]<<7)+(in_buffer[47]<<10)+(in_buffer[47]<<11))-(0-(in_buffer[48]<<2)-(in_buffer[48]<<5)+(in_buffer[48]<<8)+(in_buffer[48]<<12))-(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)+(in_buffer[49]<<7)+(in_buffer[49]<<9)+(in_buffer[49]<<12))+(0+(in_buffer[50]<<1)-(in_buffer[50]<<4)+(in_buffer[50]<<9))+(0+(in_buffer[51]<<1)+(in_buffer[51]<<3)+(in_buffer[51]<<7)+(in_buffer[51]<<10))+(0+(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<5)+(in_buffer[52]<<7)+(in_buffer[52]<<8)+(in_buffer[52]<<11)+(in_buffer[52]<<12))+(0+(in_buffer[53]<<0)+(in_buffer[53]<<6)+(in_buffer[53]<<7)+(in_buffer[53]<<11))-(0+(in_buffer[55]<<0)+(in_buffer[55]<<1)-(in_buffer[55]<<5)+(in_buffer[55]<<12))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<1)-(in_buffer[56]<<4)-(in_buffer[56]<<6)-(in_buffer[56]<<8)+(in_buffer[56]<<10)+(in_buffer[56]<<11))+(0+(in_buffer[57]<<0)+(in_buffer[57]<<1)-(in_buffer[57]<<7)+(in_buffer[57]<<9)+(in_buffer[57]<<10))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<1)-(in_buffer[58]<<4)-(in_buffer[58]<<6)-(in_buffer[58]<<8)+(in_buffer[58]<<10)+(in_buffer[58]<<11))-(0+(in_buffer[59]<<4)+(in_buffer[59]<<5)+(in_buffer[59]<<8)+(in_buffer[59]<<10))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<2)-(in_buffer[60]<<4)-(in_buffer[60]<<7)+(in_buffer[60]<<11))+(0+(in_buffer[61]<<0)+(in_buffer[61]<<4)-(in_buffer[61]<<7)+(in_buffer[61]<<10))+(0+(in_buffer[62]<<0)-(in_buffer[62]<<2)-(in_buffer[62]<<5)+(in_buffer[62]<<8)+(in_buffer[62]<<10))+(0+(in_buffer[63]<<0)-(in_buffer[63]<<2)+(in_buffer[63]<<6)-(in_buffer[63]<<8)+(in_buffer[63]<<12))-(0-(in_buffer[64]<<0)+(in_buffer[64]<<5)+(in_buffer[64]<<7)+(in_buffer[64]<<8))-(0+(in_buffer[65]<<0)+(in_buffer[65]<<1)-(in_buffer[65]<<4)-(in_buffer[65]<<6)-(in_buffer[65]<<8)+(in_buffer[65]<<10)+(in_buffer[65]<<11))-(0+(in_buffer[66]<<0)+(in_buffer[66]<<1)+(in_buffer[66]<<4)+(in_buffer[66]<<6))+(0+(in_buffer[67]<<0)+(in_buffer[67]<<2)-(in_buffer[67]<<4)-(in_buffer[67]<<7)+(in_buffer[67]<<11))+(0-(in_buffer[68]<<0)+(in_buffer[68]<<2)+(in_buffer[68]<<3)+(in_buffer[68]<<6)+(in_buffer[68]<<8)+(in_buffer[68]<<10)+(in_buffer[68]<<11))-(0+(in_buffer[69]<<0)-(in_buffer[69]<<3)+(in_buffer[69]<<8))+(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)+(in_buffer[70]<<5)+(in_buffer[70]<<11))+(0-(in_buffer[71]<<1)-(in_buffer[71]<<3)-(in_buffer[71]<<5)+(in_buffer[71]<<9)+(in_buffer[71]<<10))+(0-(in_buffer[72]<<0)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0+(in_buffer[73]<<0)+(in_buffer[73]<<3)+(in_buffer[73]<<5)+(in_buffer[73]<<9)+(in_buffer[73]<<10))+(0-(in_buffer[74]<<3)+(in_buffer[74]<<8)+(in_buffer[74]<<10)+(in_buffer[74]<<11))-(0+(in_buffer[75]<<1)+(in_buffer[75]<<4)+(in_buffer[75]<<6)+(in_buffer[75]<<10)+(in_buffer[75]<<11))+(0+(in_buffer[76]<<0)+(in_buffer[76]<<4)-(in_buffer[76]<<7)+(in_buffer[76]<<10))+(0+(in_buffer[77]<<1)-(in_buffer[77]<<3)-(in_buffer[77]<<6)+(in_buffer[77]<<9)+(in_buffer[77]<<11))-(0+(in_buffer[78]<<1)-(in_buffer[78]<<3)-(in_buffer[78]<<6)+(in_buffer[78]<<9)+(in_buffer[78]<<11))-(0-(in_buffer[79]<<0)+(in_buffer[79]<<3)-(in_buffer[79]<<5)+(in_buffer[79]<<7)+(in_buffer[79]<<8)+(in_buffer[79]<<11))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<3)+(in_buffer[80]<<6)+(in_buffer[80]<<10))+(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)+(in_buffer[81]<<7)+(in_buffer[81]<<9)+(in_buffer[81]<<12))+(0-(in_buffer[82]<<1)-(in_buffer[82]<<3)-(in_buffer[82]<<5)+(in_buffer[82]<<9)+(in_buffer[82]<<10))+(0-(in_buffer[83]<<0)+(in_buffer[83]<<4)-(in_buffer[83]<<6)-(in_buffer[83]<<8)+(in_buffer[83]<<11))-(0+(in_buffer[84]<<0)+(in_buffer[84]<<2)+(in_buffer[84]<<3)+(in_buffer[84]<<9)+(in_buffer[84]<<11))-(0+(in_buffer[85]<<0)-(in_buffer[85]<<2)-(in_buffer[85]<<5)+(in_buffer[85]<<8)+(in_buffer[85]<<10))-(0+(in_buffer[86]<<0)+(in_buffer[86]<<2)-(in_buffer[86]<<4)-(in_buffer[86]<<7)+(in_buffer[86]<<11))-(0+(in_buffer[87]<<0)+(in_buffer[87]<<3)+(in_buffer[87]<<5)+(in_buffer[87]<<9)+(in_buffer[87]<<10))+(0+(in_buffer[88]<<0)+(in_buffer[88]<<1)-(in_buffer[88]<<5)+(in_buffer[88]<<12))+(0+(in_buffer[89]<<4)+(in_buffer[89]<<5)+(in_buffer[89]<<8)+(in_buffer[89]<<10))-(0+(in_buffer[90]<<2)+(in_buffer[90]<<4)+(in_buffer[90]<<8)+(in_buffer[90]<<11))-(0+(in_buffer[91]<<0)-(in_buffer[91]<<2)-(in_buffer[91]<<5)+(in_buffer[91]<<8)+(in_buffer[91]<<10))+(0+(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<5)+(in_buffer[92]<<7)+(in_buffer[92]<<8)+(in_buffer[92]<<11)+(in_buffer[92]<<12))+(0-(in_buffer[93]<<1)+(in_buffer[93]<<4)-(in_buffer[93]<<6)+(in_buffer[93]<<8)+(in_buffer[93]<<9)+(in_buffer[93]<<12))+(0+(in_buffer[94]<<2)+(in_buffer[94]<<3)+(in_buffer[94]<<6)+(in_buffer[94]<<8))-(0-(in_buffer[95]<<0)+(in_buffer[95]<<2)+(in_buffer[95]<<3)+(in_buffer[95]<<6)+(in_buffer[95]<<8)+(in_buffer[95]<<10)+(in_buffer[95]<<11))-(0+(in_buffer[96]<<3)+(in_buffer[96]<<4)+(in_buffer[96]<<7)+(in_buffer[96]<<9))+(0+(in_buffer[97]<<4)-(in_buffer[97]<<7)+(in_buffer[97]<<12))-(0+(in_buffer[98]<<0)-(in_buffer[98]<<3)+(in_buffer[98]<<8))+(0+(in_buffer[99]<<0)+(in_buffer[99]<<2)+(in_buffer[99]<<4)-(in_buffer[99]<<6)+(in_buffer[99]<<9)+(in_buffer[99]<<12))+(0+(in_buffer[100]<<2)+(in_buffer[100]<<5)+(in_buffer[100]<<7)+(in_buffer[100]<<11)+(in_buffer[100]<<12))+(0+(in_buffer[101]<<4)+(in_buffer[101]<<5)+(in_buffer[101]<<8)+(in_buffer[101]<<10))+(0+(in_buffer[102]<<1)+(in_buffer[102]<<3)+(in_buffer[102]<<7)+(in_buffer[102]<<10))+(0+(in_buffer[103]<<0)-(in_buffer[103]<<2)+(in_buffer[103]<<5)+(in_buffer[103]<<7)+(in_buffer[103]<<8)+(in_buffer[103]<<11)+(in_buffer[103]<<12))+(0+(in_buffer[104]<<0)+(in_buffer[104]<<2)+(in_buffer[104]<<3)+(in_buffer[104]<<9)+(in_buffer[104]<<11))+(0-(in_buffer[105]<<0)-(in_buffer[105]<<2)-(in_buffer[105]<<4)+(in_buffer[105]<<8)+(in_buffer[105]<<9))-(0-(in_buffer[106]<<0)+(in_buffer[106]<<3)-(in_buffer[106]<<5)+(in_buffer[106]<<7)+(in_buffer[106]<<8)+(in_buffer[106]<<11))-(0+(in_buffer[107]<<1)+(in_buffer[107]<<7)+(in_buffer[107]<<8)+(in_buffer[107]<<12))+(0+(in_buffer[108]<<0)+(in_buffer[108]<<1)-(in_buffer[108]<<5)+(in_buffer[108]<<12))-(0+(in_buffer[109]<<2)+(in_buffer[109]<<3)+(in_buffer[109]<<6)+(in_buffer[109]<<8))-(0-(in_buffer[110]<<1)+(in_buffer[110]<<5)-(in_buffer[110]<<7)-(in_buffer[110]<<9)+(in_buffer[110]<<12))+(0-(in_buffer[111]<<0)-(in_buffer[111]<<3)+(in_buffer[111]<<6)+(in_buffer[111]<<10))+(0+(in_buffer[112]<<2)+(in_buffer[112]<<3)-(in_buffer[112]<<9)+(in_buffer[112]<<11)+(in_buffer[112]<<12))+(0+(in_buffer[113]<<0)-(in_buffer[113]<<4)-(in_buffer[113]<<9)+(in_buffer[113]<<12))-(0-(in_buffer[114]<<1)-(in_buffer[114]<<3)+(in_buffer[114]<<6)+(in_buffer[114]<<12))-(0-(in_buffer[115]<<1)+(in_buffer[115]<<3)+(in_buffer[115]<<4)+(in_buffer[115]<<7)+(in_buffer[115]<<9)+(in_buffer[115]<<11)+(in_buffer[115]<<12))-(0+(in_buffer[116]<<1)+(in_buffer[116]<<3)-(in_buffer[116]<<5)-(in_buffer[116]<<8)+(in_buffer[116]<<12))+(0-(in_buffer[118]<<2)-(in_buffer[118]<<4)-(in_buffer[118]<<6)+(in_buffer[118]<<10)+(in_buffer[118]<<11))+(0-(in_buffer[119]<<4)+(in_buffer[119]<<9)+(in_buffer[119]<<11)+(in_buffer[119]<<12))-(0-(in_buffer[120]<<0)+(in_buffer[120]<<5)+(in_buffer[120]<<7)+(in_buffer[120]<<8));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight11;
assign in_buffer_weight11=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<4)-(in_buffer[0]<<7)+(in_buffer[0]<<10))-(0-(in_buffer[1]<<0)+(in_buffer[1]<<5)+(in_buffer[1]<<7)+(in_buffer[1]<<8))-(0+(in_buffer[2]<<0)-(in_buffer[2]<<3)+(in_buffer[2]<<8))+(0+(in_buffer[4]<<0)-(in_buffer[4]<<3)+(in_buffer[4]<<8))+(0+(in_buffer[6]<<0)-(in_buffer[6]<<3)+(in_buffer[6]<<8))+(0-(in_buffer[8]<<1)+(in_buffer[8]<<6)+(in_buffer[8]<<8)+(in_buffer[8]<<9))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)+(in_buffer[9]<<6)+(in_buffer[9]<<9))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)+(in_buffer[10]<<4)+(in_buffer[10]<<6))+(0+(in_buffer[11]<<1)-(in_buffer[11]<<4)+(in_buffer[11]<<9))-(0+(in_buffer[12]<<1)-(in_buffer[12]<<4)+(in_buffer[12]<<9))+(0+(in_buffer[13]<<0)+(in_buffer[13]<<4)-(in_buffer[13]<<7)+(in_buffer[13]<<10))-(0+(in_buffer[14]<<1)+(in_buffer[14]<<2)+(in_buffer[14]<<5)+(in_buffer[14]<<7))+(0+(in_buffer[15]<<0)-(in_buffer[15]<<3)+(in_buffer[15]<<8))+(0+(in_buffer[16]<<1)-(in_buffer[16]<<4)+(in_buffer[16]<<9))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4)+(in_buffer[17]<<6))-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)-(in_buffer[18]<<4)+(in_buffer[18]<<8)+(in_buffer[18]<<9))+(0+(in_buffer[19]<<1)-(in_buffer[19]<<4)+(in_buffer[19]<<9))+(0+(in_buffer[20]<<2)+(in_buffer[20]<<3)+(in_buffer[20]<<6)+(in_buffer[20]<<8))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<1)+(in_buffer[21]<<4)+(in_buffer[21]<<6))+(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)-(in_buffer[22]<<4)+(in_buffer[22]<<8)+(in_buffer[22]<<9))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<6)+(in_buffer[23]<<9))+(0+(in_buffer[24]<<0)-(in_buffer[24]<<3)+(in_buffer[24]<<8))-(0+(in_buffer[25]<<0)+(in_buffer[25]<<2)+(in_buffer[25]<<6)+(in_buffer[25]<<9))-(0+(in_buffer[26]<<1)-(in_buffer[26]<<4)+(in_buffer[26]<<9))+(0+(in_buffer[27]<<0)+(in_buffer[27]<<2)+(in_buffer[27]<<6)+(in_buffer[27]<<9))-(0-(in_buffer[28]<<0)-(in_buffer[28]<<2)-(in_buffer[28]<<4)+(in_buffer[28]<<8)+(in_buffer[28]<<9))+(0-(in_buffer[29]<<0)+(in_buffer[29]<<5)+(in_buffer[29]<<7)+(in_buffer[29]<<8))+(0+(in_buffer[30]<<0)+(in_buffer[30]<<1)+(in_buffer[30]<<4)+(in_buffer[30]<<6))-(0+(in_buffer[31]<<2)+(in_buffer[31]<<3)+(in_buffer[31]<<6)+(in_buffer[31]<<8))-(0+(in_buffer[32]<<0)+(in_buffer[32]<<4)-(in_buffer[32]<<7)+(in_buffer[32]<<10))+(0-(in_buffer[33]<<0)-(in_buffer[33]<<2)-(in_buffer[33]<<4)+(in_buffer[33]<<8)+(in_buffer[33]<<9))-(0+(in_buffer[34]<<0)+(in_buffer[34]<<1)+(in_buffer[34]<<4)+(in_buffer[34]<<6))-(0+(in_buffer[35]<<0)+(in_buffer[35]<<4)-(in_buffer[35]<<7)+(in_buffer[35]<<10))-(0+(in_buffer[36]<<0)+(in_buffer[36]<<4)-(in_buffer[36]<<7)+(in_buffer[36]<<10))-(0+(in_buffer[37]<<0)+(in_buffer[37]<<1)+(in_buffer[37]<<4)+(in_buffer[37]<<6))-(0+(in_buffer[38]<<3)+(in_buffer[38]<<4)+(in_buffer[38]<<7)+(in_buffer[38]<<9))+(0+(in_buffer[39]<<0)+(in_buffer[39]<<1)+(in_buffer[39]<<4)+(in_buffer[39]<<6))+(0+(in_buffer[40]<<0)-(in_buffer[40]<<3)+(in_buffer[40]<<8))+(0+(in_buffer[41]<<0)+(in_buffer[41]<<1)+(in_buffer[41]<<4)+(in_buffer[41]<<6))-(0-(in_buffer[42]<<0)-(in_buffer[42]<<2)-(in_buffer[42]<<4)+(in_buffer[42]<<8)+(in_buffer[42]<<9))+(0-(in_buffer[43]<<0)+(in_buffer[43]<<5)+(in_buffer[43]<<7)+(in_buffer[43]<<8))+(0+(in_buffer[45]<<1)-(in_buffer[45]<<4)+(in_buffer[45]<<9))-(0+(in_buffer[46]<<0)+(in_buffer[46]<<1)+(in_buffer[46]<<4)+(in_buffer[46]<<6))+(0+(in_buffer[47]<<3)+(in_buffer[47]<<4)+(in_buffer[47]<<7)+(in_buffer[47]<<9))-(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)-(in_buffer[49]<<4)+(in_buffer[49]<<8)+(in_buffer[49]<<9))-(0+(in_buffer[50]<<1)-(in_buffer[50]<<4)+(in_buffer[50]<<9))-(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)-(in_buffer[51]<<4)+(in_buffer[51]<<8)+(in_buffer[51]<<9))+(0+(in_buffer[53]<<3)+(in_buffer[53]<<4)+(in_buffer[53]<<7)+(in_buffer[53]<<9))+(0+(in_buffer[54]<<0)+(in_buffer[54]<<2)+(in_buffer[54]<<6)+(in_buffer[54]<<9))-(0+(in_buffer[55]<<1)+(in_buffer[55]<<2)+(in_buffer[55]<<5)+(in_buffer[55]<<7))-(0+(in_buffer[56]<<1)-(in_buffer[56]<<4)+(in_buffer[56]<<9))+(0-(in_buffer[58]<<0)+(in_buffer[58]<<5)+(in_buffer[58]<<7)+(in_buffer[58]<<8))+(0-(in_buffer[59]<<0)+(in_buffer[59]<<5)+(in_buffer[59]<<7)+(in_buffer[59]<<8))-(0+(in_buffer[60]<<2)-(in_buffer[60]<<5)+(in_buffer[60]<<10))+(0-(in_buffer[61]<<1)+(in_buffer[61]<<6)+(in_buffer[61]<<8)+(in_buffer[61]<<9))-(0+(in_buffer[62]<<0)+(in_buffer[62]<<1)+(in_buffer[62]<<4)+(in_buffer[62]<<6))+(0+(in_buffer[63]<<3)+(in_buffer[63]<<4)+(in_buffer[63]<<7)+(in_buffer[63]<<9))+(0+(in_buffer[64]<<1)+(in_buffer[64]<<2)+(in_buffer[64]<<5)+(in_buffer[64]<<7))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)-(in_buffer[65]<<4)+(in_buffer[65]<<8)+(in_buffer[65]<<9))+(0+(in_buffer[66]<<3)+(in_buffer[66]<<4)+(in_buffer[66]<<7)+(in_buffer[66]<<9))-(0+(in_buffer[67]<<3)+(in_buffer[67]<<4)+(in_buffer[67]<<7)+(in_buffer[67]<<9))-(0+(in_buffer[68]<<1)-(in_buffer[68]<<4)+(in_buffer[68]<<9))-(0+(in_buffer[69]<<0)+(in_buffer[69]<<4)-(in_buffer[69]<<7)+(in_buffer[69]<<10))-(0+(in_buffer[70]<<1)-(in_buffer[70]<<4)+(in_buffer[70]<<9))+(0+(in_buffer[71]<<3)+(in_buffer[71]<<4)+(in_buffer[71]<<7)+(in_buffer[71]<<9))+(0-(in_buffer[72]<<0)-(in_buffer[72]<<2)-(in_buffer[72]<<4)+(in_buffer[72]<<8)+(in_buffer[72]<<9))-(0+(in_buffer[74]<<2)+(in_buffer[74]<<3)+(in_buffer[74]<<6)+(in_buffer[74]<<8))-(0+(in_buffer[75]<<2)+(in_buffer[75]<<3)+(in_buffer[75]<<6)+(in_buffer[75]<<8))+(0+(in_buffer[76]<<0)+(in_buffer[76]<<2)+(in_buffer[76]<<6)+(in_buffer[76]<<9))-(0+(in_buffer[78]<<1)+(in_buffer[78]<<2)+(in_buffer[78]<<5)+(in_buffer[78]<<7))-(0+(in_buffer[79]<<0)+(in_buffer[79]<<1)+(in_buffer[79]<<4)+(in_buffer[79]<<6))-(0+(in_buffer[80]<<0)-(in_buffer[80]<<3)+(in_buffer[80]<<8))-(0+(in_buffer[81]<<0)+(in_buffer[81]<<1)+(in_buffer[81]<<4)+(in_buffer[81]<<6))+(0-(in_buffer[82]<<0)+(in_buffer[82]<<5)+(in_buffer[82]<<7)+(in_buffer[82]<<8))-(0-(in_buffer[83]<<0)-(in_buffer[83]<<2)-(in_buffer[83]<<4)+(in_buffer[83]<<8)+(in_buffer[83]<<9))-(0+(in_buffer[84]<<1)+(in_buffer[84]<<2)+(in_buffer[84]<<5)+(in_buffer[84]<<7))-(0-(in_buffer[85]<<0)-(in_buffer[85]<<2)-(in_buffer[85]<<4)+(in_buffer[85]<<8)+(in_buffer[85]<<9))-(0+(in_buffer[86]<<0)-(in_buffer[86]<<3)+(in_buffer[86]<<8))-(0+(in_buffer[87]<<3)+(in_buffer[87]<<4)+(in_buffer[87]<<7)+(in_buffer[87]<<9))-(0+(in_buffer[88]<<0)-(in_buffer[88]<<3)+(in_buffer[88]<<8))+(0+(in_buffer[89]<<1)-(in_buffer[89]<<4)+(in_buffer[89]<<9))-(0-(in_buffer[90]<<1)+(in_buffer[90]<<6)+(in_buffer[90]<<8)+(in_buffer[90]<<9))-(0+(in_buffer[91]<<3)+(in_buffer[91]<<4)+(in_buffer[91]<<7)+(in_buffer[91]<<9))-(0-(in_buffer[92]<<1)+(in_buffer[92]<<6)+(in_buffer[92]<<8)+(in_buffer[92]<<9))+(0+(in_buffer[93]<<3)+(in_buffer[93]<<4)+(in_buffer[93]<<7)+(in_buffer[93]<<9))+(0+(in_buffer[94]<<0)+(in_buffer[94]<<2)+(in_buffer[94]<<6)+(in_buffer[94]<<9))-(0+(in_buffer[96]<<1)+(in_buffer[96]<<2)+(in_buffer[96]<<5)+(in_buffer[96]<<7))-(0+(in_buffer[97]<<2)+(in_buffer[97]<<3)+(in_buffer[97]<<6)+(in_buffer[97]<<8))-(0-(in_buffer[98]<<0)+(in_buffer[98]<<5)+(in_buffer[98]<<7)+(in_buffer[98]<<8))-(0+(in_buffer[99]<<0)+(in_buffer[99]<<2)+(in_buffer[99]<<6)+(in_buffer[99]<<9))+(0+(in_buffer[100]<<1)-(in_buffer[100]<<4)+(in_buffer[100]<<9))+(0+(in_buffer[102]<<0)-(in_buffer[102]<<3)+(in_buffer[102]<<8))+(0+(in_buffer[103]<<0)+(in_buffer[103]<<1)+(in_buffer[103]<<4)+(in_buffer[103]<<6))+(0+(in_buffer[104]<<1)+(in_buffer[104]<<2)+(in_buffer[104]<<5)+(in_buffer[104]<<7))+(0-(in_buffer[105]<<0)+(in_buffer[105]<<5)+(in_buffer[105]<<7)+(in_buffer[105]<<8))-(0+(in_buffer[106]<<0)-(in_buffer[106]<<3)+(in_buffer[106]<<8))+(0-(in_buffer[107]<<1)+(in_buffer[107]<<6)+(in_buffer[107]<<8)+(in_buffer[107]<<9))-(0+(in_buffer[109]<<2)-(in_buffer[109]<<5)+(in_buffer[109]<<10))+(0+(in_buffer[110]<<2)+(in_buffer[110]<<3)+(in_buffer[110]<<6)+(in_buffer[110]<<8))+(0-(in_buffer[111]<<1)+(in_buffer[111]<<6)+(in_buffer[111]<<8)+(in_buffer[111]<<9))+(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)-(in_buffer[112]<<4)+(in_buffer[112]<<8)+(in_buffer[112]<<9))-(0+(in_buffer[113]<<0)-(in_buffer[113]<<3)+(in_buffer[113]<<8))-(0+(in_buffer[114]<<1)-(in_buffer[114]<<4)+(in_buffer[114]<<9))-(0+(in_buffer[115]<<0)+(in_buffer[115]<<1)+(in_buffer[115]<<4)+(in_buffer[115]<<6))-(0+(in_buffer[116]<<1)-(in_buffer[116]<<4)+(in_buffer[116]<<9))+(0+(in_buffer[117]<<2)+(in_buffer[117]<<3)+(in_buffer[117]<<6)+(in_buffer[117]<<8))+(0+(in_buffer[119]<<0)+(in_buffer[119]<<1)+(in_buffer[119]<<4)+(in_buffer[119]<<6))+(0-(in_buffer[120]<<0)+(in_buffer[120]<<5)+(in_buffer[120]<<7)+(in_buffer[120]<<8));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight12;
assign in_buffer_weight12=0-(0+(in_buffer[0]<<3)+(in_buffer[0]<<5)+(in_buffer[0]<<9)+(in_buffer[0]<<12))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<1)-(in_buffer[1]<<5)+(in_buffer[1]<<12))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<2)-(in_buffer[2]<<4)-(in_buffer[2]<<6)+(in_buffer[2]<<9)+(in_buffer[2]<<10)+(in_buffer[2]<<14))+(0-(in_buffer[3]<<1)+(in_buffer[3]<<11)+(in_buffer[3]<<12))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<6)+(in_buffer[4]<<7)+(in_buffer[4]<<11))-(0+(in_buffer[5]<<2)+(in_buffer[5]<<5)+(in_buffer[5]<<7)+(in_buffer[5]<<11)+(in_buffer[5]<<12))-(0+(in_buffer[6]<<0)-(in_buffer[6]<<7)-(in_buffer[6]<<9)+(in_buffer[6]<<13))-(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)-(in_buffer[7]<<4)+(in_buffer[7]<<8)+(in_buffer[7]<<9))+(0+(in_buffer[8]<<0)-(in_buffer[8]<<4)-(in_buffer[8]<<6)+(in_buffer[8]<<8)+(in_buffer[8]<<9)+(in_buffer[8]<<13))+(0+(in_buffer[9]<<0)+(in_buffer[9]<<2)-(in_buffer[9]<<6)-(in_buffer[9]<<10)+(in_buffer[9]<<12)+(in_buffer[9]<<13))-(0-(in_buffer[10]<<1)-(in_buffer[10]<<4)+(in_buffer[10]<<7)+(in_buffer[10]<<11))+(0+(in_buffer[11]<<0)-(in_buffer[11]<<3)-(in_buffer[11]<<6)-(in_buffer[11]<<9)+(in_buffer[11]<<11)+(in_buffer[11]<<12))+(0-(in_buffer[12]<<2)-(in_buffer[12]<<4)-(in_buffer[12]<<6)+(in_buffer[12]<<10)+(in_buffer[12]<<11))+(0-(in_buffer[13]<<1)+(in_buffer[13]<<5)+(in_buffer[13]<<6)+(in_buffer[13]<<9)+(in_buffer[13]<<13))+(0+(in_buffer[14]<<5)+(in_buffer[14]<<6)+(in_buffer[14]<<9)+(in_buffer[14]<<11))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<4)-(in_buffer[15]<<6)-(in_buffer[15]<<8)+(in_buffer[15]<<11))-(0-(in_buffer[16]<<2)+(in_buffer[16]<<6)-(in_buffer[16]<<8)-(in_buffer[16]<<10)+(in_buffer[16]<<13))+(0+(in_buffer[18]<<2)+(in_buffer[18]<<4)+(in_buffer[18]<<8)+(in_buffer[18]<<11))+(0+(in_buffer[19]<<0)-(in_buffer[19]<<2)+(in_buffer[19]<<5)+(in_buffer[19]<<7)+(in_buffer[19]<<8)+(in_buffer[19]<<11)+(in_buffer[19]<<12))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<4)+(in_buffer[20]<<6)+(in_buffer[20]<<11)+(in_buffer[20]<<12))+(0-(in_buffer[21]<<0)-(in_buffer[21]<<2)-(in_buffer[21]<<10)+(in_buffer[21]<<14))-(0-(in_buffer[22]<<1)-(in_buffer[22]<<3)-(in_buffer[22]<<5)+(in_buffer[22]<<9)+(in_buffer[22]<<10))-(0-(in_buffer[23]<<0)+(in_buffer[23]<<3)+(in_buffer[23]<<5)-(in_buffer[23]<<9)+(in_buffer[23]<<13))-(0+(in_buffer[24]<<2)+(in_buffer[24]<<4)+(in_buffer[24]<<8)+(in_buffer[24]<<11))+(0+(in_buffer[25]<<4)+(in_buffer[25]<<5)+(in_buffer[25]<<8)+(in_buffer[25]<<10))-(0+(in_buffer[26]<<0)-(in_buffer[26]<<4)-(in_buffer[26]<<9)+(in_buffer[26]<<12))-(0-(in_buffer[27]<<0)+(in_buffer[27]<<3)+(in_buffer[27]<<5)-(in_buffer[27]<<9)+(in_buffer[27]<<13))-(0+(in_buffer[28]<<3)-(in_buffer[28]<<6)+(in_buffer[28]<<11))+(0+(in_buffer[29]<<5)+(in_buffer[29]<<6)+(in_buffer[29]<<9)+(in_buffer[29]<<11))+(0-(in_buffer[30]<<0)-(in_buffer[30]<<2)+(in_buffer[30]<<5)+(in_buffer[30]<<11))-(0+(in_buffer[31]<<1)+(in_buffer[31]<<5)-(in_buffer[31]<<8)+(in_buffer[31]<<11))+(0+(in_buffer[32]<<2)-(in_buffer[32]<<5)-(in_buffer[32]<<7)-(in_buffer[32]<<9)+(in_buffer[32]<<12)+(in_buffer[32]<<13))-(0-(in_buffer[33]<<0)+(in_buffer[33]<<3)-(in_buffer[33]<<6)+(in_buffer[33]<<10)+(in_buffer[33]<<12))-(0+(in_buffer[34]<<0)+(in_buffer[34]<<2)+(in_buffer[34]<<3)-(in_buffer[34]<<7)+(in_buffer[34]<<10)+(in_buffer[34]<<12)+(in_buffer[34]<<13))-(0-(in_buffer[35]<<2)-(in_buffer[35]<<5)+(in_buffer[35]<<8)+(in_buffer[35]<<12))-(0-(in_buffer[36]<<0)+(in_buffer[36]<<3)-(in_buffer[36]<<5)+(in_buffer[36]<<7)+(in_buffer[36]<<8)+(in_buffer[36]<<11))-(0+(in_buffer[37]<<1)+(in_buffer[37]<<3)-(in_buffer[37]<<5)-(in_buffer[37]<<8)+(in_buffer[37]<<12))-(0+(in_buffer[38]<<0)+(in_buffer[38]<<2)-(in_buffer[38]<<4)-(in_buffer[38]<<7)+(in_buffer[38]<<11))-(0+(in_buffer[39]<<0)+(in_buffer[39]<<1)+(in_buffer[39]<<4)+(in_buffer[39]<<6))+(0-(in_buffer[41]<<2)-(in_buffer[41]<<5)+(in_buffer[41]<<8)+(in_buffer[41]<<12))-(0+(in_buffer[42]<<0)+(in_buffer[42]<<2)-(in_buffer[42]<<5)+(in_buffer[42]<<7)+(in_buffer[42]<<8)+(in_buffer[42]<<13))+(0+(in_buffer[43]<<0)+(in_buffer[43]<<2)-(in_buffer[43]<<5)+(in_buffer[43]<<7)+(in_buffer[43]<<8)+(in_buffer[43]<<13))-(0-(in_buffer[44]<<1)-(in_buffer[44]<<3)-(in_buffer[44]<<5)+(in_buffer[44]<<9)+(in_buffer[44]<<10))-(0+(in_buffer[45]<<2)+(in_buffer[45]<<4)-(in_buffer[45]<<6)-(in_buffer[45]<<9)+(in_buffer[45]<<13))-(0+(in_buffer[46]<<3)-(in_buffer[46]<<6)+(in_buffer[46]<<11))-(0-(in_buffer[47]<<1)-(in_buffer[47]<<3)+(in_buffer[47]<<6)+(in_buffer[47]<<12))-(0+(in_buffer[48]<<0)+(in_buffer[48]<<1)+(in_buffer[48]<<4)+(in_buffer[48]<<6))+(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)-(in_buffer[49]<<4)+(in_buffer[49]<<8)+(in_buffer[49]<<9))+(0+(in_buffer[50]<<1)+(in_buffer[50]<<3)+(in_buffer[50]<<7)+(in_buffer[50]<<10))-(0-(in_buffer[51]<<0)+(in_buffer[51]<<3)+(in_buffer[51]<<4)+(in_buffer[51]<<7)-(in_buffer[51]<<9)+(in_buffer[51]<<12))+(0-(in_buffer[52]<<0)+(in_buffer[52]<<3)-(in_buffer[52]<<5)+(in_buffer[52]<<7)+(in_buffer[52]<<8)+(in_buffer[52]<<11))-(0+(in_buffer[53]<<0)+(in_buffer[53]<<1)+(in_buffer[53]<<4)+(in_buffer[53]<<8)+(in_buffer[53]<<10)+(in_buffer[53]<<12))+(0-(in_buffer[54]<<2)+(in_buffer[54]<<4)+(in_buffer[54]<<5)+(in_buffer[54]<<8)+(in_buffer[54]<<10)+(in_buffer[54]<<12)+(in_buffer[54]<<13))+(0-(in_buffer[55]<<0)+(in_buffer[55]<<3)-(in_buffer[55]<<5)+(in_buffer[55]<<7)+(in_buffer[55]<<8)+(in_buffer[55]<<11))-(0+(in_buffer[56]<<2)+(in_buffer[56]<<5)+(in_buffer[56]<<7)+(in_buffer[56]<<11)+(in_buffer[56]<<12))-(0-(in_buffer[57]<<0)-(in_buffer[57]<<3)+(in_buffer[57]<<6)+(in_buffer[57]<<10))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)-(in_buffer[58]<<4)-(in_buffer[58]<<7)+(in_buffer[58]<<11))-(0-(in_buffer[59]<<0)-(in_buffer[59]<<2)-(in_buffer[59]<<4)+(in_buffer[59]<<8)+(in_buffer[59]<<9))+(0+(in_buffer[60]<<1)+(in_buffer[60]<<2)+(in_buffer[60]<<5)+(in_buffer[60]<<7))+(0-(in_buffer[61]<<1)-(in_buffer[61]<<4)+(in_buffer[61]<<7)+(in_buffer[61]<<11))+(0-(in_buffer[62]<<3)+(in_buffer[62]<<8)+(in_buffer[62]<<10)+(in_buffer[62]<<11))+(0+(in_buffer[63]<<1)-(in_buffer[63]<<3)-(in_buffer[63]<<6)+(in_buffer[63]<<9)+(in_buffer[63]<<11))-(0+(in_buffer[64]<<0)+(in_buffer[64]<<2)+(in_buffer[64]<<6)+(in_buffer[64]<<9))+(0+(in_buffer[65]<<0)-(in_buffer[65]<<7)-(in_buffer[65]<<9)+(in_buffer[65]<<13))+(0+(in_buffer[66]<<0)-(in_buffer[66]<<3)-(in_buffer[66]<<5)-(in_buffer[66]<<7)+(in_buffer[66]<<10)+(in_buffer[66]<<11))+(0+(in_buffer[67]<<0)-(in_buffer[67]<<3)+(in_buffer[67]<<8))-(0+(in_buffer[69]<<0)+(in_buffer[69]<<1)+(in_buffer[69]<<4)+(in_buffer[69]<<6))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<4)-(in_buffer[70]<<7)+(in_buffer[70]<<10))+(0+(in_buffer[71]<<2)+(in_buffer[71]<<4)+(in_buffer[71]<<8)+(in_buffer[71]<<11))+(0-(in_buffer[72]<<0)+(in_buffer[72]<<2)+(in_buffer[72]<<3)+(in_buffer[72]<<6)+(in_buffer[72]<<8)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0-(in_buffer[73]<<1)+(in_buffer[73]<<4)-(in_buffer[73]<<6)+(in_buffer[73]<<8)+(in_buffer[73]<<9)+(in_buffer[73]<<12))+(0-(in_buffer[74]<<0)+(in_buffer[74]<<4)-(in_buffer[74]<<6)-(in_buffer[74]<<8)+(in_buffer[74]<<11))+(0+(in_buffer[75]<<2)+(in_buffer[75]<<3)+(in_buffer[75]<<6)+(in_buffer[75]<<8))+(0+(in_buffer[76]<<0)+(in_buffer[76]<<1)-(in_buffer[76]<<5)+(in_buffer[76]<<12))+(0-(in_buffer[77]<<0)+(in_buffer[77]<<4)+(in_buffer[77]<<5)+(in_buffer[77]<<8)+(in_buffer[77]<<12))+(0+(in_buffer[78]<<6)+(in_buffer[78]<<7)+(in_buffer[78]<<10)+(in_buffer[78]<<12))+(0+(in_buffer[79]<<1)-(in_buffer[79]<<3)-(in_buffer[79]<<6)+(in_buffer[79]<<9)+(in_buffer[79]<<11))-(0-(in_buffer[80]<<2)-(in_buffer[80]<<4)-(in_buffer[80]<<6)+(in_buffer[80]<<10)+(in_buffer[80]<<11))-(0+(in_buffer[81]<<1)-(in_buffer[81]<<4)+(in_buffer[81]<<9))+(0+(in_buffer[82]<<1)+(in_buffer[82]<<2)-(in_buffer[82]<<8)+(in_buffer[82]<<10)+(in_buffer[82]<<11))+(0-(in_buffer[83]<<0)+(in_buffer[83]<<10)+(in_buffer[83]<<11))+(0+(in_buffer[84]<<0)+(in_buffer[84]<<4)-(in_buffer[84]<<7)+(in_buffer[84]<<10))+(0+(in_buffer[85]<<1)+(in_buffer[85]<<5)-(in_buffer[85]<<8)+(in_buffer[85]<<11))+(0+(in_buffer[86]<<0)-(in_buffer[86]<<4)-(in_buffer[86]<<9)+(in_buffer[86]<<12))+(0+(in_buffer[87]<<0)+(in_buffer[87]<<1)+(in_buffer[87]<<5)+(in_buffer[87]<<7)+(in_buffer[87]<<10)+(in_buffer[87]<<13))+(0-(in_buffer[88]<<2)+(in_buffer[88]<<7)+(in_buffer[88]<<9)+(in_buffer[88]<<10))+(0-(in_buffer[89]<<1)+(in_buffer[89]<<5)-(in_buffer[89]<<7)-(in_buffer[89]<<9)+(in_buffer[89]<<12))-(0+(in_buffer[90]<<0)-(in_buffer[90]<<2)-(in_buffer[90]<<5)+(in_buffer[90]<<8)+(in_buffer[90]<<10))-(0+(in_buffer[91]<<0)+(in_buffer[91]<<6)+(in_buffer[91]<<7)+(in_buffer[91]<<11))+(0+(in_buffer[93]<<2)+(in_buffer[93]<<4)+(in_buffer[93]<<8)+(in_buffer[93]<<11))+(0+(in_buffer[94]<<1)+(in_buffer[94]<<2)-(in_buffer[94]<<8)+(in_buffer[94]<<10)+(in_buffer[94]<<11))-(0+(in_buffer[95]<<4)+(in_buffer[95]<<5)+(in_buffer[95]<<8)+(in_buffer[95]<<10))-(0+(in_buffer[96]<<1)-(in_buffer[96]<<3)-(in_buffer[96]<<6)+(in_buffer[96]<<9)+(in_buffer[96]<<11))+(0+(in_buffer[97]<<0)-(in_buffer[97]<<3)+(in_buffer[97]<<8))+(0-(in_buffer[98]<<0)+(in_buffer[98]<<3)-(in_buffer[98]<<5)+(in_buffer[98]<<7)+(in_buffer[98]<<8)+(in_buffer[98]<<11))-(0+(in_buffer[99]<<0)+(in_buffer[99]<<4)-(in_buffer[99]<<7)+(in_buffer[99]<<10))+(0+(in_buffer[100]<<0)+(in_buffer[100]<<2)+(in_buffer[100]<<3)+(in_buffer[100]<<9)+(in_buffer[100]<<11))+(0+(in_buffer[101]<<0)+(in_buffer[101]<<2)-(in_buffer[101]<<4)-(in_buffer[101]<<7)+(in_buffer[101]<<11))+(0+(in_buffer[102]<<0)+(in_buffer[102]<<4)-(in_buffer[102]<<7)+(in_buffer[102]<<10))+(0+(in_buffer[104]<<5)+(in_buffer[104]<<6)+(in_buffer[104]<<9)+(in_buffer[104]<<11))+(0-(in_buffer[105]<<0)-(in_buffer[105]<<3)+(in_buffer[105]<<6)+(in_buffer[105]<<10))+(0-(in_buffer[107]<<0)+(in_buffer[107]<<5)+(in_buffer[107]<<7)+(in_buffer[107]<<8))+(0+(in_buffer[108]<<0)+(in_buffer[108]<<4)-(in_buffer[108]<<7)+(in_buffer[108]<<10))+(0+(in_buffer[109]<<1)+(in_buffer[109]<<2)-(in_buffer[109]<<8)+(in_buffer[109]<<10)+(in_buffer[109]<<11))+(0+(in_buffer[110]<<0)+(in_buffer[110]<<1)+(in_buffer[110]<<4)+(in_buffer[110]<<6))+(0+(in_buffer[111]<<2)+(in_buffer[111]<<3)+(in_buffer[111]<<6)+(in_buffer[111]<<8))+(0+(in_buffer[112]<<0)-(in_buffer[112]<<4)-(in_buffer[112]<<9)+(in_buffer[112]<<12))-(0+(in_buffer[113]<<1)+(in_buffer[113]<<2)-(in_buffer[113]<<8)+(in_buffer[113]<<10)+(in_buffer[113]<<11))+(0+(in_buffer[114]<<0)+(in_buffer[114]<<1)-(in_buffer[114]<<4)-(in_buffer[114]<<6)-(in_buffer[114]<<8)+(in_buffer[114]<<10)+(in_buffer[114]<<11))+(0+(in_buffer[115]<<0)-(in_buffer[115]<<2)+(in_buffer[115]<<5)+(in_buffer[115]<<7)+(in_buffer[115]<<8)+(in_buffer[115]<<11)+(in_buffer[115]<<12))-(0+(in_buffer[116]<<2)+(in_buffer[116]<<3)+(in_buffer[116]<<6)+(in_buffer[116]<<8))-(0+(in_buffer[117]<<4)+(in_buffer[117]<<5)+(in_buffer[117]<<8)+(in_buffer[117]<<10))+(0+(in_buffer[118]<<1)+(in_buffer[118]<<4)+(in_buffer[118]<<6)+(in_buffer[118]<<10)+(in_buffer[118]<<11))-(0-(in_buffer[119]<<0)+(in_buffer[119]<<3)+(in_buffer[119]<<4)+(in_buffer[119]<<7)-(in_buffer[119]<<9)+(in_buffer[119]<<12))+(0+(in_buffer[120]<<0)-(in_buffer[120]<<3)+(in_buffer[120]<<8));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight13;
assign in_buffer_weight13=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3)-(in_buffer[0]<<7)+(in_buffer[0]<<10)+(in_buffer[0]<<12)+(in_buffer[0]<<13))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<6)+(in_buffer[1]<<9)+(in_buffer[1]<<10)+(in_buffer[1]<<13))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<6)+(in_buffer[2]<<7)+(in_buffer[2]<<11))+(0-(in_buffer[3]<<2)+(in_buffer[3]<<12)+(in_buffer[3]<<13))+(0+(in_buffer[4]<<0)-(in_buffer[4]<<4)-(in_buffer[4]<<9)+(in_buffer[4]<<12))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<5)+(in_buffer[5]<<7)+(in_buffer[5]<<10)+(in_buffer[5]<<11))+(0+(in_buffer[6]<<0)-(in_buffer[6]<<4)-(in_buffer[6]<<9)+(in_buffer[6]<<12))+(0-(in_buffer[7]<<1)+(in_buffer[7]<<4)-(in_buffer[7]<<6)+(in_buffer[7]<<8)+(in_buffer[7]<<9)+(in_buffer[7]<<12))+(0-(in_buffer[8]<<2)+(in_buffer[8]<<7)+(in_buffer[8]<<9)+(in_buffer[8]<<10))-(0+(in_buffer[9]<<1)+(in_buffer[9]<<5)-(in_buffer[9]<<8)+(in_buffer[9]<<11))-(0+(in_buffer[10]<<2)+(in_buffer[10]<<4)+(in_buffer[10]<<8)+(in_buffer[10]<<11))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<6)+(in_buffer[11]<<8)+(in_buffer[11]<<10)+(in_buffer[11]<<13))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<3)-(in_buffer[12]<<6)-(in_buffer[12]<<8)+(in_buffer[12]<<13))+(0-(in_buffer[13]<<0)+(in_buffer[13]<<3)-(in_buffer[13]<<5)+(in_buffer[13]<<7)+(in_buffer[13]<<8)+(in_buffer[13]<<11))+(0+(in_buffer[14]<<2)+(in_buffer[14]<<3)+(in_buffer[14]<<6)+(in_buffer[14]<<8))-(0+(in_buffer[15]<<0)-(in_buffer[15]<<3)-(in_buffer[15]<<5)-(in_buffer[15]<<7)+(in_buffer[15]<<10)+(in_buffer[15]<<11))+(0+(in_buffer[16]<<1)-(in_buffer[16]<<4)+(in_buffer[16]<<9))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)-(in_buffer[17]<<7)+(in_buffer[17]<<9)+(in_buffer[17]<<10))-(0+(in_buffer[18]<<3)-(in_buffer[18]<<6)+(in_buffer[18]<<11))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<5)+(in_buffer[19]<<7)+(in_buffer[19]<<8))+(0+(in_buffer[20]<<4)-(in_buffer[20]<<7)+(in_buffer[20]<<12))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<6)+(in_buffer[21]<<8)+(in_buffer[21]<<10)+(in_buffer[21]<<13))-(0+(in_buffer[22]<<1)+(in_buffer[22]<<2)-(in_buffer[22]<<5)-(in_buffer[22]<<7)-(in_buffer[22]<<9)+(in_buffer[22]<<11)+(in_buffer[22]<<12))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<2)-(in_buffer[23]<<5)-(in_buffer[23]<<7)-(in_buffer[23]<<9)+(in_buffer[23]<<11)+(in_buffer[23]<<12))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<10)+(in_buffer[24]<<11))+(0+(in_buffer[25]<<4)-(in_buffer[25]<<7)+(in_buffer[25]<<12))-(0-(in_buffer[26]<<0)+(in_buffer[26]<<10)+(in_buffer[26]<<11))-(0-(in_buffer[27]<<0)-(in_buffer[27]<<3)+(in_buffer[27]<<6)+(in_buffer[27]<<10))-(0-(in_buffer[28]<<2)-(in_buffer[28]<<4)-(in_buffer[28]<<6)+(in_buffer[28]<<10)+(in_buffer[28]<<11))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<3)+(in_buffer[29]<<7)+(in_buffer[29]<<12))+(0+(in_buffer[30]<<0)+(in_buffer[30]<<2)-(in_buffer[30]<<4)-(in_buffer[30]<<7)+(in_buffer[30]<<11))+(0-(in_buffer[31]<<1)-(in_buffer[31]<<3)-(in_buffer[31]<<5)+(in_buffer[31]<<9)+(in_buffer[31]<<10))-(0+(in_buffer[32]<<2)-(in_buffer[32]<<4)-(in_buffer[32]<<7)+(in_buffer[32]<<10)+(in_buffer[32]<<12))-(0+(in_buffer[33]<<3)-(in_buffer[33]<<6)+(in_buffer[33]<<11))+(0-(in_buffer[34]<<0)-(in_buffer[34]<<3)+(in_buffer[34]<<8)+(in_buffer[34]<<11)+(in_buffer[34]<<12))+(0+(in_buffer[35]<<0)-(in_buffer[35]<<2)+(in_buffer[35]<<5)+(in_buffer[35]<<7)+(in_buffer[35]<<8)+(in_buffer[35]<<11)+(in_buffer[35]<<12))+(0+(in_buffer[36]<<1)+(in_buffer[36]<<7)+(in_buffer[36]<<8)+(in_buffer[36]<<12))-(0-(in_buffer[37]<<1)-(in_buffer[37]<<3)+(in_buffer[37]<<8)+(in_buffer[37]<<10)+(in_buffer[37]<<13))-(0+(in_buffer[38]<<0)-(in_buffer[38]<<4)-(in_buffer[38]<<9)+(in_buffer[38]<<12))-(0+(in_buffer[39]<<0)-(in_buffer[39]<<3)-(in_buffer[39]<<5)-(in_buffer[39]<<7)+(in_buffer[39]<<10)+(in_buffer[39]<<11))+(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)-(in_buffer[40]<<4)+(in_buffer[40]<<8)+(in_buffer[40]<<9))+(0+(in_buffer[41]<<0)-(in_buffer[41]<<2)-(in_buffer[41]<<4)+(in_buffer[41]<<7)+(in_buffer[41]<<10)+(in_buffer[41]<<12))+(0+(in_buffer[42]<<2)+(in_buffer[42]<<4)+(in_buffer[42]<<8)+(in_buffer[42]<<11))-(0+(in_buffer[43]<<0)-(in_buffer[43]<<3)-(in_buffer[43]<<6)-(in_buffer[43]<<9)+(in_buffer[43]<<11)+(in_buffer[43]<<12))+(0-(in_buffer[44]<<2)+(in_buffer[44]<<7)+(in_buffer[44]<<9)+(in_buffer[44]<<10))+(0-(in_buffer[45]<<0)+(in_buffer[45]<<4)-(in_buffer[45]<<7)-(in_buffer[45]<<10)+(in_buffer[45]<<13))-(0+(in_buffer[46]<<0)+(in_buffer[46]<<2)+(in_buffer[46]<<6)+(in_buffer[46]<<9))-(0+(in_buffer[47]<<0)-(in_buffer[47]<<2)-(in_buffer[47]<<5)+(in_buffer[47]<<8)+(in_buffer[47]<<10))-(0+(in_buffer[48]<<3)+(in_buffer[48]<<7)-(in_buffer[48]<<10)+(in_buffer[48]<<13))-(0+(in_buffer[49]<<2)-(in_buffer[49]<<5)+(in_buffer[49]<<10))-(0+(in_buffer[50]<<3)-(in_buffer[50]<<6)+(in_buffer[50]<<11))-(0+(in_buffer[51]<<2)+(in_buffer[51]<<4)+(in_buffer[51]<<8)+(in_buffer[51]<<11))+(0-(in_buffer[52]<<0)+(in_buffer[52]<<3)+(in_buffer[52]<<5)-(in_buffer[52]<<9)+(in_buffer[52]<<13))+(0+(in_buffer[53]<<1)-(in_buffer[53]<<3)-(in_buffer[53]<<6)+(in_buffer[53]<<9)+(in_buffer[53]<<11))-(0-(in_buffer[54]<<1)+(in_buffer[54]<<3)+(in_buffer[54]<<4)+(in_buffer[54]<<7)+(in_buffer[54]<<9)+(in_buffer[54]<<11)+(in_buffer[54]<<12))-(0-(in_buffer[55]<<0)+(in_buffer[55]<<5)-(in_buffer[55]<<8)-(in_buffer[55]<<10)+(in_buffer[55]<<12)+(in_buffer[55]<<13))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<3)+(in_buffer[56]<<9)+(in_buffer[56]<<11))-(0+(in_buffer[57]<<3)-(in_buffer[57]<<5)-(in_buffer[57]<<8)+(in_buffer[57]<<11)+(in_buffer[57]<<13))-(0-(in_buffer[58]<<0)+(in_buffer[58]<<3)+(in_buffer[58]<<4)+(in_buffer[58]<<7)-(in_buffer[58]<<9)+(in_buffer[58]<<12))-(0+(in_buffer[59]<<3)+(in_buffer[59]<<4)+(in_buffer[59]<<7)+(in_buffer[59]<<9))+(0+(in_buffer[60]<<0)+(in_buffer[60]<<3)+(in_buffer[60]<<5)+(in_buffer[60]<<9)+(in_buffer[60]<<10))+(0+(in_buffer[61]<<0)+(in_buffer[61]<<2)-(in_buffer[61]<<4)-(in_buffer[61]<<7)+(in_buffer[61]<<11))-(0+(in_buffer[62]<<0)+(in_buffer[62]<<1)-(in_buffer[62]<<7)+(in_buffer[62]<<9)+(in_buffer[62]<<10))+(0+(in_buffer[63]<<0)+(in_buffer[63]<<2)+(in_buffer[63]<<6)+(in_buffer[63]<<9))+(0+(in_buffer[64]<<0)+(in_buffer[64]<<3)+(in_buffer[64]<<5)+(in_buffer[64]<<9)+(in_buffer[64]<<10))+(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)-(in_buffer[65]<<4)+(in_buffer[65]<<8)+(in_buffer[65]<<9))-(0+(in_buffer[66]<<3)+(in_buffer[66]<<5)+(in_buffer[66]<<9)+(in_buffer[66]<<12))+(0-(in_buffer[67]<<0)+(in_buffer[67]<<5)+(in_buffer[67]<<6)-(in_buffer[67]<<9)+(in_buffer[67]<<11)+(in_buffer[67]<<12))-(0-(in_buffer[68]<<0)-(in_buffer[68]<<2)-(in_buffer[68]<<5)+(in_buffer[68]<<8)-(in_buffer[68]<<10)+(in_buffer[68]<<13))+(0-(in_buffer[69]<<1)-(in_buffer[69]<<3)-(in_buffer[69]<<5)+(in_buffer[69]<<9)+(in_buffer[69]<<10))+(0-(in_buffer[70]<<1)+(in_buffer[70]<<11)+(in_buffer[70]<<12))+(0+(in_buffer[71]<<1)+(in_buffer[71]<<4)+(in_buffer[71]<<6)+(in_buffer[71]<<10)+(in_buffer[71]<<11))+(0-(in_buffer[72]<<3)+(in_buffer[72]<<8)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0-(in_buffer[73]<<0)-(in_buffer[73]<<3)+(in_buffer[73]<<6)+(in_buffer[73]<<10))+(0-(in_buffer[74]<<0)+(in_buffer[74]<<5)+(in_buffer[74]<<7)+(in_buffer[74]<<8))+(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)-(in_buffer[75]<<4)+(in_buffer[75]<<8)+(in_buffer[75]<<9))+(0+(in_buffer[76]<<1)+(in_buffer[76]<<2)+(in_buffer[76]<<5)+(in_buffer[76]<<7))-(0+(in_buffer[77]<<1)+(in_buffer[77]<<2)+(in_buffer[77]<<5)+(in_buffer[77]<<7))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<2)-(in_buffer[78]<<4)-(in_buffer[78]<<6)+(in_buffer[78]<<11)+(in_buffer[78]<<12))-(0-(in_buffer[79]<<1)-(in_buffer[79]<<3)+(in_buffer[79]<<6)+(in_buffer[79]<<12))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<3)+(in_buffer[80]<<8)+(in_buffer[80]<<11)+(in_buffer[80]<<12))+(0+(in_buffer[81]<<1)+(in_buffer[81]<<3)+(in_buffer[81]<<4)+(in_buffer[81]<<10)+(in_buffer[81]<<12))-(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<5)+(in_buffer[82]<<11))+(0+(in_buffer[83]<<1)+(in_buffer[83]<<2)+(in_buffer[83]<<5)+(in_buffer[83]<<7))-(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)-(in_buffer[84]<<4)+(in_buffer[84]<<8)+(in_buffer[84]<<9))-(0+(in_buffer[85]<<3)+(in_buffer[85]<<4)+(in_buffer[85]<<7)+(in_buffer[85]<<9))+(0+(in_buffer[86]<<0)+(in_buffer[86]<<4)-(in_buffer[86]<<7)+(in_buffer[86]<<10))-(0-(in_buffer[87]<<1)+(in_buffer[87]<<6)+(in_buffer[87]<<8)+(in_buffer[87]<<9))+(0-(in_buffer[88]<<2)-(in_buffer[88]<<5)+(in_buffer[88]<<8)+(in_buffer[88]<<12))+(0-(in_buffer[89]<<0)+(in_buffer[89]<<4)-(in_buffer[89]<<6)-(in_buffer[89]<<8)+(in_buffer[89]<<11))-(0+(in_buffer[90]<<0)+(in_buffer[90]<<2)-(in_buffer[90]<<5)+(in_buffer[90]<<7)+(in_buffer[90]<<8)+(in_buffer[90]<<13))+(0-(in_buffer[91]<<0)+(in_buffer[91]<<4)-(in_buffer[91]<<6)-(in_buffer[91]<<8)+(in_buffer[91]<<11))+(0+(in_buffer[92]<<0)+(in_buffer[92]<<4)+(in_buffer[92]<<6)+(in_buffer[92]<<11)+(in_buffer[92]<<12))-(0-(in_buffer[94]<<0)+(in_buffer[94]<<5)+(in_buffer[94]<<7)+(in_buffer[94]<<8))+(0-(in_buffer[95]<<1)+(in_buffer[95]<<4)-(in_buffer[95]<<6)+(in_buffer[95]<<8)+(in_buffer[95]<<9)+(in_buffer[95]<<12))-(0+(in_buffer[96]<<0)+(in_buffer[96]<<1)-(in_buffer[96]<<7)+(in_buffer[96]<<9)+(in_buffer[96]<<10))+(0-(in_buffer[97]<<0)+(in_buffer[97]<<4)-(in_buffer[97]<<6)-(in_buffer[97]<<8)+(in_buffer[97]<<11))+(0-(in_buffer[98]<<2)-(in_buffer[98]<<4)-(in_buffer[98]<<6)+(in_buffer[98]<<10)+(in_buffer[98]<<11))+(0+(in_buffer[99]<<0)+(in_buffer[99]<<2)+(in_buffer[99]<<3)-(in_buffer[99]<<6)-(in_buffer[99]<<8)+(in_buffer[99]<<13))-(0-(in_buffer[100]<<1)+(in_buffer[100]<<6)+(in_buffer[100]<<8)+(in_buffer[100]<<9))-(0+(in_buffer[101]<<1)+(in_buffer[101]<<3)+(in_buffer[101]<<7)+(in_buffer[101]<<10))+(0-(in_buffer[102]<<0)+(in_buffer[102]<<4)-(in_buffer[102]<<6)-(in_buffer[102]<<8)+(in_buffer[102]<<11))+(0-(in_buffer[103]<<0)+(in_buffer[103]<<5)+(in_buffer[103]<<6)-(in_buffer[103]<<9)+(in_buffer[103]<<11)+(in_buffer[103]<<12))+(0+(in_buffer[104]<<1)-(in_buffer[104]<<3)-(in_buffer[104]<<6)+(in_buffer[104]<<9)+(in_buffer[104]<<11))+(0+(in_buffer[105]<<0)+(in_buffer[105]<<2)+(in_buffer[105]<<6)+(in_buffer[105]<<9))+(0-(in_buffer[106]<<2)-(in_buffer[106]<<4)-(in_buffer[106]<<6)+(in_buffer[106]<<10)+(in_buffer[106]<<11))-(0-(in_buffer[107]<<1)+(in_buffer[107]<<6)+(in_buffer[107]<<8)+(in_buffer[107]<<9))-(0+(in_buffer[108]<<1)-(in_buffer[108]<<3)-(in_buffer[108]<<6)+(in_buffer[108]<<9)+(in_buffer[108]<<11))+(0+(in_buffer[109]<<0)-(in_buffer[109]<<3)-(in_buffer[109]<<6)-(in_buffer[109]<<9)+(in_buffer[109]<<11)+(in_buffer[109]<<12))+(0+(in_buffer[110]<<0)+(in_buffer[110]<<1)-(in_buffer[110]<<5)+(in_buffer[110]<<12))-(0+(in_buffer[111]<<1)+(in_buffer[111]<<4)+(in_buffer[111]<<8)+(in_buffer[111]<<13))-(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)+(in_buffer[112]<<5)+(in_buffer[112]<<11))-(0+(in_buffer[113]<<3)+(in_buffer[113]<<5)+(in_buffer[113]<<9)+(in_buffer[113]<<12))+(0+(in_buffer[114]<<0)+(in_buffer[114]<<2)-(in_buffer[114]<<4)-(in_buffer[114]<<7)+(in_buffer[114]<<11))+(0-(in_buffer[115]<<0)+(in_buffer[115]<<6)+(in_buffer[115]<<7)+(in_buffer[115]<<13))+(0+(in_buffer[116]<<1)+(in_buffer[116]<<6)+(in_buffer[116]<<9)+(in_buffer[116]<<10)+(in_buffer[116]<<13))+(0+(in_buffer[117]<<1)+(in_buffer[117]<<2)-(in_buffer[117]<<5)-(in_buffer[117]<<7)-(in_buffer[117]<<9)+(in_buffer[117]<<11)+(in_buffer[117]<<12))+(0+(in_buffer[118]<<1)-(in_buffer[118]<<4)-(in_buffer[118]<<6)-(in_buffer[118]<<8)+(in_buffer[118]<<11)+(in_buffer[118]<<12))+(0+(in_buffer[119]<<0)+(in_buffer[119]<<3)+(in_buffer[119]<<7)+(in_buffer[119]<<12))+(0+(in_buffer[120]<<0)+(in_buffer[120]<<2)-(in_buffer[120]<<4)+(in_buffer[120]<<8)+(in_buffer[120]<<12)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight14;
assign in_buffer_weight14=0-(0-(in_buffer[0]<<0)-(in_buffer[0]<<4)+(in_buffer[0]<<9)+(in_buffer[0]<<10)+(in_buffer[0]<<13))+(0-(in_buffer[1]<<0)+(in_buffer[1]<<4)-(in_buffer[1]<<6)-(in_buffer[1]<<8)+(in_buffer[1]<<11))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<1)-(in_buffer[2]<<4)-(in_buffer[2]<<6)-(in_buffer[2]<<8)+(in_buffer[2]<<10)+(in_buffer[2]<<11))-(0-(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<7)+(in_buffer[3]<<9)+(in_buffer[3]<<12))-(0+(in_buffer[4]<<1)+(in_buffer[4]<<3)-(in_buffer[4]<<5)-(in_buffer[4]<<8)+(in_buffer[4]<<12))+(0+(in_buffer[5]<<1)-(in_buffer[5]<<3)+(in_buffer[5]<<7)-(in_buffer[5]<<9)+(in_buffer[5]<<13))-(0+(in_buffer[6]<<1)+(in_buffer[6]<<2)-(in_buffer[6]<<5)-(in_buffer[6]<<7)-(in_buffer[6]<<9)+(in_buffer[6]<<11)+(in_buffer[6]<<12))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<3)+(in_buffer[7]<<6)+(in_buffer[7]<<8)+(in_buffer[7]<<10)+(in_buffer[7]<<13))-(0+(in_buffer[8]<<0)+(in_buffer[8]<<2)+(in_buffer[8]<<4)-(in_buffer[8]<<6)+(in_buffer[8]<<9)+(in_buffer[8]<<12))+(0+(in_buffer[9]<<2)+(in_buffer[9]<<4)-(in_buffer[9]<<6)-(in_buffer[9]<<9)+(in_buffer[9]<<13))+(0-(in_buffer[10]<<1)+(in_buffer[10]<<4)-(in_buffer[10]<<7)+(in_buffer[10]<<11)+(in_buffer[10]<<13))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<5)-(in_buffer[11]<<9)+(in_buffer[11]<<13))-(0-(in_buffer[12]<<0)-(in_buffer[12]<<2)-(in_buffer[12]<<4)-(in_buffer[12]<<6)+(in_buffer[12]<<11)+(in_buffer[12]<<12))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<4)-(in_buffer[13]<<6)-(in_buffer[13]<<8)+(in_buffer[13]<<11))+(0-(in_buffer[14]<<3)+(in_buffer[14]<<8)+(in_buffer[14]<<10)+(in_buffer[14]<<11))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<4)-(in_buffer[15]<<6)-(in_buffer[15]<<8)+(in_buffer[15]<<11))+(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<3)+(in_buffer[16]<<9)+(in_buffer[16]<<11))-(0+(in_buffer[17]<<2)-(in_buffer[17]<<5)+(in_buffer[17]<<10))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<5)-(in_buffer[18]<<7)-(in_buffer[18]<<9)+(in_buffer[18]<<12))-(0+(in_buffer[19]<<2)+(in_buffer[19]<<4)+(in_buffer[19]<<8)+(in_buffer[19]<<11))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<7)-(in_buffer[20]<<9)+(in_buffer[20]<<13))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<1)-(in_buffer[21]<<5)+(in_buffer[21]<<8)+(in_buffer[21]<<9)+(in_buffer[21]<<13)+(in_buffer[21]<<14))-(0-(in_buffer[22]<<0)-(in_buffer[22]<<3)+(in_buffer[22]<<6)+(in_buffer[22]<<10))-(0+(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<7)+(in_buffer[23]<<8)+(in_buffer[23]<<11)+(in_buffer[23]<<12))-(0+(in_buffer[24]<<1)-(in_buffer[24]<<5)-(in_buffer[24]<<10)+(in_buffer[24]<<13))-(0+(in_buffer[25]<<0)-(in_buffer[25]<<4)-(in_buffer[25]<<9)+(in_buffer[25]<<12))-(0-(in_buffer[27]<<0)+(in_buffer[27]<<4)-(in_buffer[27]<<6)-(in_buffer[27]<<8)+(in_buffer[27]<<11))-(0+(in_buffer[28]<<0)+(in_buffer[28]<<2)+(in_buffer[28]<<6)+(in_buffer[28]<<9))-(0+(in_buffer[29]<<1)-(in_buffer[29]<<3)-(in_buffer[29]<<6)+(in_buffer[29]<<9)+(in_buffer[29]<<11))-(0-(in_buffer[30]<<1)-(in_buffer[30]<<4)+(in_buffer[30]<<7)+(in_buffer[30]<<11))-(0-(in_buffer[31]<<0)+(in_buffer[31]<<10)+(in_buffer[31]<<11))+(0-(in_buffer[32]<<1)+(in_buffer[32]<<7)+(in_buffer[32]<<8)+(in_buffer[32]<<14))-(0+(in_buffer[33]<<0)+(in_buffer[33]<<2)+(in_buffer[33]<<3)+(in_buffer[33]<<9)+(in_buffer[33]<<11))-(0-(in_buffer[34]<<0)+(in_buffer[34]<<3)-(in_buffer[34]<<6)+(in_buffer[34]<<10)+(in_buffer[34]<<12))-(0-(in_buffer[35]<<1)-(in_buffer[35]<<3)+(in_buffer[35]<<6)+(in_buffer[35]<<12))-(0+(in_buffer[36]<<1)+(in_buffer[36]<<3)+(in_buffer[36]<<7)+(in_buffer[36]<<10))-(0+(in_buffer[37]<<0)-(in_buffer[37]<<4)-(in_buffer[37]<<9)+(in_buffer[37]<<12))-(0-(in_buffer[38]<<1)-(in_buffer[38]<<3)-(in_buffer[38]<<5)+(in_buffer[38]<<9)+(in_buffer[38]<<10))-(0-(in_buffer[39]<<0)+(in_buffer[39]<<3)-(in_buffer[39]<<5)+(in_buffer[39]<<7)+(in_buffer[39]<<8)+(in_buffer[39]<<11))-(0+(in_buffer[40]<<1)+(in_buffer[40]<<2)+(in_buffer[40]<<5)+(in_buffer[40]<<7))+(0+(in_buffer[41]<<0)-(in_buffer[41]<<3)+(in_buffer[41]<<8))+(0-(in_buffer[42]<<2)-(in_buffer[42]<<4)-(in_buffer[42]<<6)+(in_buffer[42]<<10)+(in_buffer[42]<<11))+(0-(in_buffer[43]<<0)-(in_buffer[43]<<2)-(in_buffer[43]<<4)+(in_buffer[43]<<7)-(in_buffer[43]<<10)+(in_buffer[43]<<12)+(in_buffer[43]<<13))-(0-(in_buffer[44]<<1)-(in_buffer[44]<<3)-(in_buffer[44]<<5)+(in_buffer[44]<<9)+(in_buffer[44]<<10))-(0-(in_buffer[45]<<3)+(in_buffer[45]<<8)+(in_buffer[45]<<10)+(in_buffer[45]<<11))+(0+(in_buffer[46]<<1)+(in_buffer[46]<<2)+(in_buffer[46]<<5)+(in_buffer[46]<<7))+(0+(in_buffer[47]<<2)+(in_buffer[47]<<4)+(in_buffer[47]<<8)+(in_buffer[47]<<11))-(0+(in_buffer[48]<<0)+(in_buffer[48]<<3)+(in_buffer[48]<<5)+(in_buffer[48]<<9)+(in_buffer[48]<<10))+(0+(in_buffer[49]<<0)+(in_buffer[49]<<3)+(in_buffer[49]<<5)+(in_buffer[49]<<9)+(in_buffer[49]<<10))-(0-(in_buffer[50]<<0)-(in_buffer[50]<<3)+(in_buffer[50]<<6)+(in_buffer[50]<<10))+(0+(in_buffer[51]<<0)+(in_buffer[51]<<6)+(in_buffer[51]<<7)+(in_buffer[51]<<11))-(0-(in_buffer[52]<<0)+(in_buffer[52]<<5)+(in_buffer[52]<<7)+(in_buffer[52]<<8))+(0+(in_buffer[53]<<0)+(in_buffer[53]<<1)+(in_buffer[53]<<4)+(in_buffer[53]<<6))+(0+(in_buffer[54]<<1)+(in_buffer[54]<<3)+(in_buffer[54]<<6)+(in_buffer[54]<<8)+(in_buffer[54]<<11)+(in_buffer[54]<<12))-(0-(in_buffer[55]<<1)+(in_buffer[55]<<5)-(in_buffer[55]<<7)-(in_buffer[55]<<9)+(in_buffer[55]<<12))-(0+(in_buffer[56]<<0)-(in_buffer[56]<<4)-(in_buffer[56]<<9)+(in_buffer[56]<<12))+(0-(in_buffer[57]<<0)+(in_buffer[57]<<5)+(in_buffer[57]<<7)+(in_buffer[57]<<8))+(0+(in_buffer[58]<<0)-(in_buffer[58]<<2)+(in_buffer[58]<<6)-(in_buffer[58]<<8)+(in_buffer[58]<<12))+(0+(in_buffer[59]<<0)+(in_buffer[59]<<3)+(in_buffer[59]<<5)+(in_buffer[59]<<9)+(in_buffer[59]<<10))+(0+(in_buffer[60]<<1)+(in_buffer[60]<<3)-(in_buffer[60]<<5)-(in_buffer[60]<<8)+(in_buffer[60]<<12))-(0+(in_buffer[61]<<0)+(in_buffer[61]<<2)-(in_buffer[61]<<4)-(in_buffer[61]<<7)+(in_buffer[61]<<11))+(0-(in_buffer[62]<<1)+(in_buffer[62]<<3)+(in_buffer[62]<<4)+(in_buffer[62]<<7)+(in_buffer[62]<<9)+(in_buffer[62]<<11)+(in_buffer[62]<<12))-(0+(in_buffer[63]<<0)-(in_buffer[63]<<3)+(in_buffer[63]<<8))-(0+(in_buffer[65]<<0)-(in_buffer[65]<<2)-(in_buffer[65]<<5)+(in_buffer[65]<<8)+(in_buffer[65]<<10))+(0+(in_buffer[66]<<0)+(in_buffer[66]<<6)+(in_buffer[66]<<7)+(in_buffer[66]<<11))+(0+(in_buffer[67]<<1)-(in_buffer[67]<<3)-(in_buffer[67]<<6)+(in_buffer[67]<<9)+(in_buffer[67]<<11))-(0-(in_buffer[68]<<0)+(in_buffer[68]<<5)+(in_buffer[68]<<7)+(in_buffer[68]<<8))+(0+(in_buffer[69]<<3)-(in_buffer[69]<<6)+(in_buffer[69]<<11))+(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)-(in_buffer[70]<<4)+(in_buffer[70]<<8)+(in_buffer[70]<<9))+(0+(in_buffer[71]<<5)+(in_buffer[71]<<6)+(in_buffer[71]<<9)+(in_buffer[71]<<11))-(0-(in_buffer[72]<<1)+(in_buffer[72]<<6)+(in_buffer[72]<<8)+(in_buffer[72]<<9))+(0+(in_buffer[73]<<2)+(in_buffer[73]<<3)-(in_buffer[73]<<9)+(in_buffer[73]<<11)+(in_buffer[73]<<12))-(0+(in_buffer[74]<<0)-(in_buffer[74]<<3)+(in_buffer[74]<<8))+(0-(in_buffer[75]<<0)+(in_buffer[75]<<3)-(in_buffer[75]<<5)+(in_buffer[75]<<7)+(in_buffer[75]<<8)+(in_buffer[75]<<11))+(0-(in_buffer[77]<<0)+(in_buffer[77]<<5)+(in_buffer[77]<<7)+(in_buffer[77]<<8))+(0+(in_buffer[78]<<0)-(in_buffer[78]<<2)+(in_buffer[78]<<6)-(in_buffer[78]<<8)+(in_buffer[78]<<12))-(0+(in_buffer[79]<<2)+(in_buffer[79]<<3)+(in_buffer[79]<<6)+(in_buffer[79]<<8))+(0+(in_buffer[80]<<0)+(in_buffer[80]<<6)+(in_buffer[80]<<7)+(in_buffer[80]<<11))+(0+(in_buffer[81]<<0)-(in_buffer[81]<<2)-(in_buffer[81]<<5)+(in_buffer[81]<<8)+(in_buffer[81]<<10))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)-(in_buffer[82]<<4)-(in_buffer[82]<<6)+(in_buffer[82]<<11)+(in_buffer[82]<<12))+(0+(in_buffer[83]<<0)+(in_buffer[83]<<1)+(in_buffer[83]<<4)+(in_buffer[83]<<6))+(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)+(in_buffer[84]<<7)+(in_buffer[84]<<9)+(in_buffer[84]<<12))-(0+(in_buffer[85]<<1)+(in_buffer[85]<<2)+(in_buffer[85]<<5)+(in_buffer[85]<<7))+(0+(in_buffer[86]<<0)-(in_buffer[86]<<3)-(in_buffer[86]<<5)-(in_buffer[86]<<7)+(in_buffer[86]<<10)+(in_buffer[86]<<11))+(0+(in_buffer[87]<<2)+(in_buffer[87]<<4)+(in_buffer[87]<<8)+(in_buffer[87]<<11))-(0-(in_buffer[88]<<0)+(in_buffer[88]<<3)-(in_buffer[88]<<6)+(in_buffer[88]<<10)+(in_buffer[88]<<12))+(0+(in_buffer[89]<<0)+(in_buffer[89]<<1)+(in_buffer[89]<<4)+(in_buffer[89]<<6))+(0+(in_buffer[90]<<1)+(in_buffer[90]<<2)+(in_buffer[90]<<5)+(in_buffer[90]<<7))+(0-(in_buffer[91]<<0)+(in_buffer[91]<<3)+(in_buffer[91]<<4)+(in_buffer[91]<<7)-(in_buffer[91]<<9)+(in_buffer[91]<<12))-(0+(in_buffer[92]<<2)+(in_buffer[92]<<3)+(in_buffer[92]<<6)+(in_buffer[92]<<8))+(0-(in_buffer[93]<<3)+(in_buffer[93]<<8)+(in_buffer[93]<<10)+(in_buffer[93]<<11))-(0-(in_buffer[94]<<0)-(in_buffer[94]<<2)+(in_buffer[94]<<5)+(in_buffer[94]<<11))-(0+(in_buffer[95]<<0)+(in_buffer[95]<<4)-(in_buffer[95]<<7)+(in_buffer[95]<<10))-(0+(in_buffer[96]<<0)-(in_buffer[96]<<2)-(in_buffer[96]<<5)+(in_buffer[96]<<8)+(in_buffer[96]<<10))+(0+(in_buffer[97]<<1)-(in_buffer[97]<<4)+(in_buffer[97]<<9))+(0-(in_buffer[98]<<0)+(in_buffer[98]<<5)+(in_buffer[98]<<7)+(in_buffer[98]<<8))-(0-(in_buffer[99]<<0)+(in_buffer[99]<<3)-(in_buffer[99]<<5)+(in_buffer[99]<<7)+(in_buffer[99]<<8)+(in_buffer[99]<<11))+(0-(in_buffer[101]<<2)-(in_buffer[101]<<4)-(in_buffer[101]<<6)+(in_buffer[101]<<10)+(in_buffer[101]<<11))+(0+(in_buffer[102]<<0)+(in_buffer[102]<<3)+(in_buffer[102]<<7)+(in_buffer[102]<<12))-(0+(in_buffer[103]<<0)+(in_buffer[103]<<6)+(in_buffer[103]<<7)+(in_buffer[103]<<11))+(0+(in_buffer[104]<<2)+(in_buffer[104]<<3)+(in_buffer[104]<<6)+(in_buffer[104]<<8))-(0+(in_buffer[105]<<1)+(in_buffer[105]<<4)+(in_buffer[105]<<6)+(in_buffer[105]<<10)+(in_buffer[105]<<11))+(0+(in_buffer[106]<<3)+(in_buffer[106]<<4)+(in_buffer[106]<<7)+(in_buffer[106]<<9))+(0+(in_buffer[107]<<0)+(in_buffer[107]<<3)+(in_buffer[107]<<5)+(in_buffer[107]<<9)+(in_buffer[107]<<10))+(0-(in_buffer[108]<<2)+(in_buffer[108]<<7)+(in_buffer[108]<<9)+(in_buffer[108]<<10))-(0+(in_buffer[109]<<2)+(in_buffer[109]<<6)-(in_buffer[109]<<9)+(in_buffer[109]<<12))+(0-(in_buffer[110]<<0)-(in_buffer[110]<<3)+(in_buffer[110]<<6)+(in_buffer[110]<<10))+(0+(in_buffer[111]<<0)+(in_buffer[111]<<1)-(in_buffer[111]<<5)+(in_buffer[111]<<12))+(0+(in_buffer[112]<<0)-(in_buffer[112]<<3)+(in_buffer[112]<<8))-(0-(in_buffer[113]<<0)+(in_buffer[113]<<3)-(in_buffer[113]<<5)+(in_buffer[113]<<7)+(in_buffer[113]<<8)+(in_buffer[113]<<11))+(0-(in_buffer[114]<<0)+(in_buffer[114]<<10)+(in_buffer[114]<<11))+(0-(in_buffer[115]<<4)+(in_buffer[115]<<9)+(in_buffer[115]<<11)+(in_buffer[115]<<12))-(0-(in_buffer[116]<<1)-(in_buffer[116]<<3)+(in_buffer[116]<<6)+(in_buffer[116]<<12))-(0+(in_buffer[117]<<0)-(in_buffer[117]<<2)-(in_buffer[117]<<4)+(in_buffer[117]<<7)+(in_buffer[117]<<10)+(in_buffer[117]<<12))-(0-(in_buffer[118]<<0)-(in_buffer[118]<<3)+(in_buffer[118]<<8)+(in_buffer[118]<<11)+(in_buffer[118]<<12))-(0+(in_buffer[119]<<0)+(in_buffer[119]<<2)+(in_buffer[119]<<3)+(in_buffer[119]<<9)+(in_buffer[119]<<11))-(0-(in_buffer[120]<<1)+(in_buffer[120]<<3)+(in_buffer[120]<<4)+(in_buffer[120]<<7)+(in_buffer[120]<<9)+(in_buffer[120]<<11)+(in_buffer[120]<<12));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight15;
assign in_buffer_weight15=0-(0+(in_buffer[0]<<3)+(in_buffer[0]<<7)-(in_buffer[0]<<10)+(in_buffer[0]<<13))+(0+(in_buffer[1]<<1)+(in_buffer[1]<<3)+(in_buffer[1]<<4)+(in_buffer[1]<<10)+(in_buffer[1]<<12))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<3)+(in_buffer[2]<<6)+(in_buffer[2]<<8)+(in_buffer[2]<<11)+(in_buffer[2]<<12))+(0-(in_buffer[3]<<1)+(in_buffer[3]<<5)-(in_buffer[3]<<7)-(in_buffer[3]<<9)+(in_buffer[3]<<12))+(0+(in_buffer[4]<<2)+(in_buffer[4]<<4)+(in_buffer[4]<<8)+(in_buffer[4]<<11))+(0+(in_buffer[5]<<0)-(in_buffer[5]<<4)-(in_buffer[5]<<9)+(in_buffer[5]<<12))-(0-(in_buffer[6]<<0)+(in_buffer[6]<<10)+(in_buffer[6]<<11))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<2)+(in_buffer[7]<<6)+(in_buffer[7]<<9))+(0+(in_buffer[8]<<1)+(in_buffer[8]<<2)+(in_buffer[8]<<5)+(in_buffer[8]<<7))+(0+(in_buffer[9]<<3)+(in_buffer[9]<<4)+(in_buffer[9]<<7)+(in_buffer[9]<<9))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<4)+(in_buffer[10]<<8)+(in_buffer[10]<<13))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<7)+(in_buffer[11]<<9)+(in_buffer[11]<<12))-(0-(in_buffer[12]<<0)-(in_buffer[12]<<3)+(in_buffer[12]<<8)+(in_buffer[12]<<11)+(in_buffer[12]<<12))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2)-(in_buffer[13]<<4)-(in_buffer[13]<<7)+(in_buffer[13]<<11))+(0-(in_buffer[14]<<0)+(in_buffer[14]<<4)-(in_buffer[14]<<7)-(in_buffer[14]<<10)+(in_buffer[14]<<13))+(0+(in_buffer[15]<<0)-(in_buffer[15]<<4)-(in_buffer[15]<<9)+(in_buffer[15]<<12))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<5)+(in_buffer[16]<<7)+(in_buffer[16]<<8))+(0-(in_buffer[17]<<0)+(in_buffer[17]<<5)+(in_buffer[17]<<7)+(in_buffer[17]<<8))-(0+(in_buffer[18]<<0)-(in_buffer[18]<<3)+(in_buffer[18]<<8))-(0+(in_buffer[19]<<0)-(in_buffer[19]<<2)-(in_buffer[19]<<4)+(in_buffer[19]<<7)+(in_buffer[19]<<10)+(in_buffer[19]<<12))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<3)+(in_buffer[20]<<4)+(in_buffer[20]<<7)+(in_buffer[20]<<8)+(in_buffer[20]<<11)+(in_buffer[20]<<14))-(0-(in_buffer[21]<<0)+(in_buffer[21]<<4)-(in_buffer[21]<<6)-(in_buffer[21]<<8)+(in_buffer[21]<<11))-(0-(in_buffer[22]<<0)+(in_buffer[22]<<4)+(in_buffer[22]<<5)+(in_buffer[22]<<8)+(in_buffer[22]<<12))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<7)+(in_buffer[23]<<10)+(in_buffer[23]<<11))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<10)+(in_buffer[24]<<11))+(0-(in_buffer[25]<<0)+(in_buffer[25]<<5)+(in_buffer[25]<<6)-(in_buffer[25]<<9)+(in_buffer[25]<<11)+(in_buffer[25]<<12))+(0+(in_buffer[26]<<1)+(in_buffer[26]<<3)+(in_buffer[26]<<5)-(in_buffer[26]<<7)+(in_buffer[26]<<10)+(in_buffer[26]<<13))+(0-(in_buffer[27]<<0)+(in_buffer[27]<<3)+(in_buffer[27]<<4)+(in_buffer[27]<<7)-(in_buffer[27]<<9)+(in_buffer[27]<<12))-(0+(in_buffer[28]<<2)+(in_buffer[28]<<3)+(in_buffer[28]<<6)+(in_buffer[28]<<8))-(0-(in_buffer[29]<<1)+(in_buffer[29]<<4)+(in_buffer[29]<<5)+(in_buffer[29]<<8)-(in_buffer[29]<<10)+(in_buffer[29]<<13))-(0+(in_buffer[30]<<4)+(in_buffer[30]<<5)+(in_buffer[30]<<8)+(in_buffer[30]<<10))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<1)+(in_buffer[31]<<4)-(in_buffer[31]<<6)+(in_buffer[31]<<9)+(in_buffer[31]<<11)+(in_buffer[31]<<13))-(0-(in_buffer[32]<<2)-(in_buffer[32]<<4)+(in_buffer[32]<<7)+(in_buffer[32]<<13))+(0+(in_buffer[33]<<2)+(in_buffer[33]<<4)+(in_buffer[33]<<8)+(in_buffer[33]<<11))+(0+(in_buffer[34]<<0)-(in_buffer[34]<<3)+(in_buffer[34]<<8))+(0+(in_buffer[35]<<2)+(in_buffer[35]<<4)+(in_buffer[35]<<8)+(in_buffer[35]<<11))+(0-(in_buffer[36]<<1)-(in_buffer[36]<<3)-(in_buffer[36]<<5)+(in_buffer[36]<<9)+(in_buffer[36]<<10))+(0-(in_buffer[37]<<0)+(in_buffer[37]<<5)+(in_buffer[37]<<6)-(in_buffer[37]<<9)+(in_buffer[37]<<11)+(in_buffer[37]<<12))+(0+(in_buffer[38]<<0)+(in_buffer[38]<<1)-(in_buffer[38]<<5)+(in_buffer[38]<<12))-(0-(in_buffer[39]<<0)+(in_buffer[39]<<4)+(in_buffer[39]<<5)+(in_buffer[39]<<8)+(in_buffer[39]<<12))-(0+(in_buffer[40]<<0)+(in_buffer[40]<<4)+(in_buffer[40]<<6)+(in_buffer[40]<<11)+(in_buffer[40]<<12))+(0-(in_buffer[41]<<1)-(in_buffer[41]<<3)-(in_buffer[41]<<5)+(in_buffer[41]<<9)+(in_buffer[41]<<10))-(0-(in_buffer[42]<<0)+(in_buffer[42]<<10)+(in_buffer[42]<<11))-(0+(in_buffer[43]<<0)+(in_buffer[43]<<3)+(in_buffer[43]<<5)+(in_buffer[43]<<9)+(in_buffer[43]<<10))+(0+(in_buffer[44]<<0)-(in_buffer[44]<<7)-(in_buffer[44]<<9)+(in_buffer[44]<<13))+(0-(in_buffer[45]<<0)-(in_buffer[45]<<2)+(in_buffer[45]<<7)+(in_buffer[45]<<9)+(in_buffer[45]<<12))+(0-(in_buffer[46]<<0)+(in_buffer[46]<<2)+(in_buffer[46]<<3)+(in_buffer[46]<<9)+(in_buffer[46]<<13))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<4)-(in_buffer[47]<<7)+(in_buffer[47]<<10))+(0+(in_buffer[49]<<0)-(in_buffer[49]<<4)-(in_buffer[49]<<9)+(in_buffer[49]<<12))-(0-(in_buffer[50]<<0)-(in_buffer[50]<<3)+(in_buffer[50]<<6)+(in_buffer[50]<<10))-(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)+(in_buffer[51]<<5)+(in_buffer[51]<<11))+(0+(in_buffer[52]<<0)-(in_buffer[52]<<3)-(in_buffer[52]<<6)-(in_buffer[52]<<9)+(in_buffer[52]<<11)+(in_buffer[52]<<12))-(0+(in_buffer[53]<<1)+(in_buffer[53]<<5)-(in_buffer[53]<<8)+(in_buffer[53]<<11))-(0+(in_buffer[54]<<1)+(in_buffer[54]<<2)+(in_buffer[54]<<5)+(in_buffer[54]<<7))-(0+(in_buffer[55]<<1)+(in_buffer[55]<<3)+(in_buffer[55]<<4)+(in_buffer[55]<<10)+(in_buffer[55]<<12))+(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<6)+(in_buffer[56]<<9))+(0+(in_buffer[57]<<3)+(in_buffer[57]<<5)+(in_buffer[57]<<9)+(in_buffer[57]<<12))+(0+(in_buffer[58]<<1)+(in_buffer[58]<<3)+(in_buffer[58]<<7)+(in_buffer[58]<<10))+(0+(in_buffer[59]<<2)-(in_buffer[59]<<5)+(in_buffer[59]<<10))+(0+(in_buffer[60]<<0)-(in_buffer[60]<<4)-(in_buffer[60]<<9)+(in_buffer[60]<<12))-(0+(in_buffer[61]<<0)+(in_buffer[61]<<3)+(in_buffer[61]<<5)+(in_buffer[61]<<9)+(in_buffer[61]<<10))+(0+(in_buffer[62]<<1)+(in_buffer[62]<<3)+(in_buffer[62]<<7)+(in_buffer[62]<<10))+(0+(in_buffer[63]<<2)+(in_buffer[63]<<6)-(in_buffer[63]<<9)+(in_buffer[63]<<12))-(0+(in_buffer[64]<<3)-(in_buffer[64]<<6)+(in_buffer[64]<<11))-(0+(in_buffer[65]<<0)-(in_buffer[65]<<3)-(in_buffer[65]<<5)-(in_buffer[65]<<7)+(in_buffer[65]<<10)+(in_buffer[65]<<11))-(0-(in_buffer[66]<<1)+(in_buffer[66]<<4)-(in_buffer[66]<<6)+(in_buffer[66]<<8)+(in_buffer[66]<<9)+(in_buffer[66]<<12))+(0+(in_buffer[67]<<0)+(in_buffer[67]<<6)+(in_buffer[67]<<7)+(in_buffer[67]<<11))+(0-(in_buffer[68]<<0)+(in_buffer[68]<<3)-(in_buffer[68]<<5)+(in_buffer[68]<<7)+(in_buffer[68]<<8)+(in_buffer[68]<<11))+(0-(in_buffer[69]<<0)-(in_buffer[69]<<3)+(in_buffer[69]<<6)+(in_buffer[69]<<10))-(0-(in_buffer[70]<<0)-(in_buffer[70]<<3)+(in_buffer[70]<<6)+(in_buffer[70]<<10))+(0+(in_buffer[71]<<0)+(in_buffer[71]<<1)-(in_buffer[71]<<7)+(in_buffer[71]<<9)+(in_buffer[71]<<10))-(0-(in_buffer[72]<<0)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0+(in_buffer[73]<<2)+(in_buffer[73]<<3)+(in_buffer[73]<<6)+(in_buffer[73]<<8))+(0-(in_buffer[74]<<3)+(in_buffer[74]<<8)+(in_buffer[74]<<10)+(in_buffer[74]<<11))-(0-(in_buffer[75]<<0)+(in_buffer[75]<<10)+(in_buffer[75]<<11))+(0+(in_buffer[76]<<0)+(in_buffer[76]<<4)-(in_buffer[76]<<7)+(in_buffer[76]<<10))-(0-(in_buffer[77]<<0)-(in_buffer[77]<<2)-(in_buffer[77]<<4)+(in_buffer[77]<<8)+(in_buffer[77]<<9))+(0+(in_buffer[78]<<5)+(in_buffer[78]<<6)+(in_buffer[78]<<9)+(in_buffer[78]<<11))+(0-(in_buffer[79]<<3)-(in_buffer[79]<<5)-(in_buffer[79]<<7)+(in_buffer[79]<<11)+(in_buffer[79]<<12))+(0-(in_buffer[80]<<0)+(in_buffer[80]<<5)+(in_buffer[80]<<7)+(in_buffer[80]<<8))+(0+(in_buffer[81]<<1)+(in_buffer[81]<<5)-(in_buffer[81]<<8)+(in_buffer[81]<<11))+(0+(in_buffer[82]<<4)-(in_buffer[82]<<7)+(in_buffer[82]<<12))+(0-(in_buffer[83]<<2)+(in_buffer[83]<<7)+(in_buffer[83]<<9)+(in_buffer[83]<<10))+(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)+(in_buffer[84]<<5)+(in_buffer[84]<<11))+(0+(in_buffer[85]<<5)-(in_buffer[85]<<8)+(in_buffer[85]<<13))+(0+(in_buffer[86]<<0)-(in_buffer[86]<<3)-(in_buffer[86]<<5)-(in_buffer[86]<<7)+(in_buffer[86]<<10)+(in_buffer[86]<<11))-(0+(in_buffer[87]<<0)-(in_buffer[87]<<2)-(in_buffer[87]<<5)+(in_buffer[87]<<8)+(in_buffer[87]<<10))-(0-(in_buffer[88]<<0)-(in_buffer[88]<<3)+(in_buffer[88]<<6)+(in_buffer[88]<<10))-(0-(in_buffer[89]<<1)-(in_buffer[89]<<3)-(in_buffer[89]<<5)+(in_buffer[89]<<9)+(in_buffer[89]<<10))+(0+(in_buffer[90]<<0)+(in_buffer[90]<<2)-(in_buffer[90]<<8)+(in_buffer[90]<<11)+(in_buffer[90]<<12))-(0+(in_buffer[91]<<1)+(in_buffer[91]<<3)+(in_buffer[91]<<7)+(in_buffer[91]<<10))+(0+(in_buffer[92]<<0)+(in_buffer[92]<<4)-(in_buffer[92]<<7)+(in_buffer[92]<<10))-(0+(in_buffer[93]<<0)-(in_buffer[93]<<3)+(in_buffer[93]<<8))-(0-(in_buffer[94]<<0)+(in_buffer[94]<<3)+(in_buffer[94]<<4)+(in_buffer[94]<<7)-(in_buffer[94]<<9)+(in_buffer[94]<<12))-(0+(in_buffer[95]<<0)+(in_buffer[95]<<4)-(in_buffer[95]<<7)+(in_buffer[95]<<10))+(0-(in_buffer[96]<<0)+(in_buffer[96]<<6)+(in_buffer[96]<<7)+(in_buffer[96]<<13))+(0+(in_buffer[97]<<3)+(in_buffer[97]<<5)+(in_buffer[97]<<9)+(in_buffer[97]<<12))+(0+(in_buffer[98]<<1)+(in_buffer[98]<<3)+(in_buffer[98]<<7)+(in_buffer[98]<<10))-(0+(in_buffer[99]<<0)-(in_buffer[99]<<2)+(in_buffer[99]<<5)+(in_buffer[99]<<7)+(in_buffer[99]<<8)+(in_buffer[99]<<11)+(in_buffer[99]<<12))+(0-(in_buffer[100]<<3)+(in_buffer[100]<<8)+(in_buffer[100]<<10)+(in_buffer[100]<<11))+(0+(in_buffer[101]<<0)+(in_buffer[101]<<2)-(in_buffer[101]<<4)+(in_buffer[101]<<8)+(in_buffer[101]<<12)+(in_buffer[101]<<13))+(0-(in_buffer[102]<<0)-(in_buffer[102]<<3)+(in_buffer[102]<<6)+(in_buffer[102]<<10))-(0+(in_buffer[103]<<0)-(in_buffer[103]<<2)-(in_buffer[103]<<5)+(in_buffer[103]<<8)+(in_buffer[103]<<10))-(0-(in_buffer[104]<<2)+(in_buffer[104]<<7)+(in_buffer[104]<<9)+(in_buffer[104]<<10))+(0-(in_buffer[105]<<1)+(in_buffer[105]<<6)+(in_buffer[105]<<8)+(in_buffer[105]<<9))+(0+(in_buffer[106]<<0)+(in_buffer[106]<<6)+(in_buffer[106]<<7)+(in_buffer[106]<<11))+(0+(in_buffer[107]<<1)+(in_buffer[107]<<3)+(in_buffer[107]<<5)-(in_buffer[107]<<7)+(in_buffer[107]<<10)+(in_buffer[107]<<13))+(0+(in_buffer[108]<<2)+(in_buffer[108]<<6)-(in_buffer[108]<<9)+(in_buffer[108]<<12))-(0+(in_buffer[109]<<2)+(in_buffer[109]<<6)-(in_buffer[109]<<9)+(in_buffer[109]<<12))-(0+(in_buffer[110]<<0)+(in_buffer[110]<<5)+(in_buffer[110]<<8)+(in_buffer[110]<<9)+(in_buffer[110]<<12))+(0+(in_buffer[111]<<1)-(in_buffer[111]<<4)+(in_buffer[111]<<9))+(0+(in_buffer[112]<<3)+(in_buffer[112]<<7)-(in_buffer[112]<<10)+(in_buffer[112]<<13))-(0-(in_buffer[113]<<1)+(in_buffer[113]<<6)+(in_buffer[113]<<8)+(in_buffer[113]<<9))+(0+(in_buffer[114]<<0)+(in_buffer[114]<<2)+(in_buffer[114]<<6)+(in_buffer[114]<<9))-(0+(in_buffer[115]<<4)+(in_buffer[115]<<5)+(in_buffer[115]<<8)+(in_buffer[115]<<10))+(0-(in_buffer[116]<<0)-(in_buffer[116]<<2)+(in_buffer[116]<<5)+(in_buffer[116]<<11))-(0+(in_buffer[117]<<1)+(in_buffer[117]<<2)+(in_buffer[117]<<5)+(in_buffer[117]<<7))-(0-(in_buffer[119]<<0)-(in_buffer[119]<<2)-(in_buffer[119]<<4)+(in_buffer[119]<<8)+(in_buffer[119]<<9))-(0+(in_buffer[120]<<2)+(in_buffer[120]<<3)-(in_buffer[120]<<9)+(in_buffer[120]<<11)+(in_buffer[120]<<12));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight16;
assign in_buffer_weight16=0-(0+(in_buffer[0]<<1)+(in_buffer[0]<<2)+(in_buffer[0]<<5)+(in_buffer[0]<<7))-(0-(in_buffer[1]<<1)+(in_buffer[1]<<6)+(in_buffer[1]<<8)+(in_buffer[1]<<9))-(0-(in_buffer[2]<<0)+(in_buffer[2]<<5)+(in_buffer[2]<<7)+(in_buffer[2]<<8))+(0+(in_buffer[3]<<3)+(in_buffer[3]<<4)+(in_buffer[3]<<7)+(in_buffer[3]<<9))-(0+(in_buffer[4]<<0)-(in_buffer[4]<<3)+(in_buffer[4]<<8))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<2)+(in_buffer[5]<<5)+(in_buffer[5]<<7))+(0+(in_buffer[6]<<1)-(in_buffer[6]<<4)+(in_buffer[6]<<9))-(0+(in_buffer[7]<<2)+(in_buffer[7]<<3)+(in_buffer[7]<<6)+(in_buffer[7]<<8))-(0-(in_buffer[8]<<0)-(in_buffer[8]<<2)-(in_buffer[8]<<4)+(in_buffer[8]<<8)+(in_buffer[8]<<9))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<1)+(in_buffer[9]<<4)+(in_buffer[9]<<6))-(0-(in_buffer[10]<<0)-(in_buffer[10]<<2)-(in_buffer[10]<<4)+(in_buffer[10]<<8)+(in_buffer[10]<<9))+(0-(in_buffer[11]<<0)-(in_buffer[11]<<2)-(in_buffer[11]<<4)+(in_buffer[11]<<8)+(in_buffer[11]<<9))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<2)+(in_buffer[12]<<6)+(in_buffer[12]<<9))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<3)+(in_buffer[14]<<6)+(in_buffer[14]<<8))-(0-(in_buffer[15]<<0)+(in_buffer[15]<<5)+(in_buffer[15]<<7)+(in_buffer[15]<<8))+(0+(in_buffer[16]<<3)+(in_buffer[16]<<4)+(in_buffer[16]<<7)+(in_buffer[16]<<9))-(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)-(in_buffer[17]<<4)+(in_buffer[17]<<8)+(in_buffer[17]<<9))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<2)+(in_buffer[19]<<6)+(in_buffer[19]<<9))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<3)+(in_buffer[20]<<8))-(0+(in_buffer[21]<<0)-(in_buffer[21]<<3)+(in_buffer[21]<<8))-(0+(in_buffer[22]<<1)-(in_buffer[22]<<4)+(in_buffer[22]<<9))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<7))-(0-(in_buffer[24]<<0)+(in_buffer[24]<<5)+(in_buffer[24]<<7)+(in_buffer[24]<<8))+(0+(in_buffer[25]<<3)+(in_buffer[25]<<4)+(in_buffer[25]<<7)+(in_buffer[25]<<9))-(0-(in_buffer[26]<<0)+(in_buffer[26]<<5)+(in_buffer[26]<<7)+(in_buffer[26]<<8))-(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)-(in_buffer[27]<<4)+(in_buffer[27]<<8)+(in_buffer[27]<<9))-(0+(in_buffer[28]<<1)-(in_buffer[28]<<4)+(in_buffer[28]<<9))-(0-(in_buffer[29]<<1)+(in_buffer[29]<<6)+(in_buffer[29]<<8)+(in_buffer[29]<<9))-(0+(in_buffer[30]<<0)+(in_buffer[30]<<4)-(in_buffer[30]<<7)+(in_buffer[30]<<10))-(0+(in_buffer[31]<<0)-(in_buffer[31]<<3)+(in_buffer[31]<<8))+(0+(in_buffer[32]<<2)+(in_buffer[32]<<3)+(in_buffer[32]<<6)+(in_buffer[32]<<8))+(0+(in_buffer[33]<<1)+(in_buffer[33]<<2)+(in_buffer[33]<<5)+(in_buffer[33]<<7))+(0-(in_buffer[34]<<0)-(in_buffer[34]<<2)-(in_buffer[34]<<4)+(in_buffer[34]<<8)+(in_buffer[34]<<9))+(0+(in_buffer[35]<<2)+(in_buffer[35]<<3)+(in_buffer[35]<<6)+(in_buffer[35]<<8))-(0+(in_buffer[36]<<1)+(in_buffer[36]<<2)+(in_buffer[36]<<5)+(in_buffer[36]<<7))-(0-(in_buffer[37]<<0)-(in_buffer[37]<<2)-(in_buffer[37]<<4)+(in_buffer[37]<<8)+(in_buffer[37]<<9))+(0-(in_buffer[38]<<0)-(in_buffer[38]<<2)-(in_buffer[38]<<4)+(in_buffer[38]<<8)+(in_buffer[38]<<9))-(0+(in_buffer[39]<<2)-(in_buffer[39]<<5)+(in_buffer[39]<<10))+(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)-(in_buffer[40]<<4)+(in_buffer[40]<<8)+(in_buffer[40]<<9))-(0-(in_buffer[41]<<1)+(in_buffer[41]<<6)+(in_buffer[41]<<8)+(in_buffer[41]<<9))+(0+(in_buffer[43]<<0)+(in_buffer[43]<<1)+(in_buffer[43]<<4)+(in_buffer[43]<<6))-(0+(in_buffer[44]<<1)-(in_buffer[44]<<4)+(in_buffer[44]<<9))+(0-(in_buffer[46]<<1)+(in_buffer[46]<<6)+(in_buffer[46]<<8)+(in_buffer[46]<<9))-(0+(in_buffer[47]<<2)+(in_buffer[47]<<3)+(in_buffer[47]<<6)+(in_buffer[47]<<8))-(0+(in_buffer[48]<<2)+(in_buffer[48]<<3)+(in_buffer[48]<<6)+(in_buffer[48]<<8))-(0+(in_buffer[49]<<1)+(in_buffer[49]<<2)+(in_buffer[49]<<5)+(in_buffer[49]<<7))+(0+(in_buffer[50]<<1)+(in_buffer[50]<<2)+(in_buffer[50]<<5)+(in_buffer[50]<<7))-(0+(in_buffer[51]<<0)+(in_buffer[51]<<1)+(in_buffer[51]<<4)+(in_buffer[51]<<6))+(0+(in_buffer[52]<<2)+(in_buffer[52]<<3)+(in_buffer[52]<<6)+(in_buffer[52]<<8))+(0+(in_buffer[54]<<0)+(in_buffer[54]<<2)+(in_buffer[54]<<6)+(in_buffer[54]<<9))+(0+(in_buffer[55]<<0)+(in_buffer[55]<<2)+(in_buffer[55]<<6)+(in_buffer[55]<<9))-(0+(in_buffer[56]<<1)-(in_buffer[56]<<4)+(in_buffer[56]<<9))-(0+(in_buffer[57]<<2)+(in_buffer[57]<<3)+(in_buffer[57]<<6)+(in_buffer[57]<<8))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)+(in_buffer[58]<<6)+(in_buffer[58]<<9))-(0-(in_buffer[59]<<0)-(in_buffer[59]<<2)-(in_buffer[59]<<4)+(in_buffer[59]<<8)+(in_buffer[59]<<9))+(0+(in_buffer[60]<<0)-(in_buffer[60]<<3)+(in_buffer[60]<<8))+(0+(in_buffer[61]<<1)-(in_buffer[61]<<4)+(in_buffer[61]<<9))+(0+(in_buffer[62]<<1)-(in_buffer[62]<<4)+(in_buffer[62]<<9))+(0-(in_buffer[64]<<0)+(in_buffer[64]<<5)+(in_buffer[64]<<7)+(in_buffer[64]<<8))-(0-(in_buffer[65]<<0)-(in_buffer[65]<<2)-(in_buffer[65]<<4)+(in_buffer[65]<<8)+(in_buffer[65]<<9))-(0-(in_buffer[66]<<0)+(in_buffer[66]<<5)+(in_buffer[66]<<7)+(in_buffer[66]<<8))+(0-(in_buffer[67]<<0)-(in_buffer[67]<<2)-(in_buffer[67]<<4)+(in_buffer[67]<<8)+(in_buffer[67]<<9))+(0-(in_buffer[68]<<0)+(in_buffer[68]<<5)+(in_buffer[68]<<7)+(in_buffer[68]<<8))+(0-(in_buffer[69]<<0)+(in_buffer[69]<<5)+(in_buffer[69]<<7)+(in_buffer[69]<<8))-(0+(in_buffer[71]<<0)-(in_buffer[71]<<3)+(in_buffer[71]<<8))-(0+(in_buffer[72]<<0)+(in_buffer[72]<<1)+(in_buffer[72]<<4)+(in_buffer[72]<<6))-(0+(in_buffer[73]<<0)+(in_buffer[73]<<4)-(in_buffer[73]<<7)+(in_buffer[73]<<10))+(0-(in_buffer[74]<<0)+(in_buffer[74]<<5)+(in_buffer[74]<<7)+(in_buffer[74]<<8))-(0-(in_buffer[75]<<0)-(in_buffer[75]<<2)-(in_buffer[75]<<4)+(in_buffer[75]<<8)+(in_buffer[75]<<9))+(0+(in_buffer[76]<<2)+(in_buffer[76]<<3)+(in_buffer[76]<<6)+(in_buffer[76]<<8))-(0+(in_buffer[77]<<0)+(in_buffer[77]<<1)+(in_buffer[77]<<4)+(in_buffer[77]<<6))-(0-(in_buffer[78]<<1)+(in_buffer[78]<<6)+(in_buffer[78]<<8)+(in_buffer[78]<<9))+(0+(in_buffer[79]<<1)-(in_buffer[79]<<4)+(in_buffer[79]<<9))-(0+(in_buffer[80]<<1)-(in_buffer[80]<<4)+(in_buffer[80]<<9))+(0+(in_buffer[81]<<0)+(in_buffer[81]<<2)+(in_buffer[81]<<6)+(in_buffer[81]<<9))-(0+(in_buffer[82]<<1)+(in_buffer[82]<<2)+(in_buffer[82]<<5)+(in_buffer[82]<<7))-(0-(in_buffer[83]<<0)+(in_buffer[83]<<5)+(in_buffer[83]<<7)+(in_buffer[83]<<8))-(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)-(in_buffer[84]<<4)+(in_buffer[84]<<8)+(in_buffer[84]<<9))-(0+(in_buffer[85]<<0)+(in_buffer[85]<<2)+(in_buffer[85]<<6)+(in_buffer[85]<<9))+(0-(in_buffer[87]<<0)-(in_buffer[87]<<2)-(in_buffer[87]<<4)+(in_buffer[87]<<8)+(in_buffer[87]<<9))-(0-(in_buffer[88]<<0)-(in_buffer[88]<<2)-(in_buffer[88]<<4)+(in_buffer[88]<<8)+(in_buffer[88]<<9))-(0+(in_buffer[89]<<1)-(in_buffer[89]<<4)+(in_buffer[89]<<9))-(0+(in_buffer[90]<<2)+(in_buffer[90]<<3)+(in_buffer[90]<<6)+(in_buffer[90]<<8))+(0-(in_buffer[91]<<0)-(in_buffer[91]<<2)-(in_buffer[91]<<4)+(in_buffer[91]<<8)+(in_buffer[91]<<9))+(0-(in_buffer[92]<<1)+(in_buffer[92]<<6)+(in_buffer[92]<<8)+(in_buffer[92]<<9))-(0+(in_buffer[93]<<0)+(in_buffer[93]<<4)-(in_buffer[93]<<7)+(in_buffer[93]<<10))+(0+(in_buffer[94]<<1)-(in_buffer[94]<<4)+(in_buffer[94]<<9))+(0+(in_buffer[95]<<1)+(in_buffer[95]<<2)+(in_buffer[95]<<5)+(in_buffer[95]<<7))+(0+(in_buffer[96]<<2)+(in_buffer[96]<<3)+(in_buffer[96]<<6)+(in_buffer[96]<<8))-(0+(in_buffer[97]<<1)-(in_buffer[97]<<4)+(in_buffer[97]<<9))-(0+(in_buffer[98]<<1)-(in_buffer[98]<<4)+(in_buffer[98]<<9))+(0+(in_buffer[99]<<2)+(in_buffer[99]<<3)+(in_buffer[99]<<6)+(in_buffer[99]<<8))-(0-(in_buffer[101]<<1)+(in_buffer[101]<<6)+(in_buffer[101]<<8)+(in_buffer[101]<<9))-(0-(in_buffer[102]<<0)+(in_buffer[102]<<5)+(in_buffer[102]<<7)+(in_buffer[102]<<8))+(0+(in_buffer[104]<<1)-(in_buffer[104]<<4)+(in_buffer[104]<<9))-(0+(in_buffer[105]<<3)+(in_buffer[105]<<4)+(in_buffer[105]<<7)+(in_buffer[105]<<9))-(0+(in_buffer[106]<<3)+(in_buffer[106]<<4)+(in_buffer[106]<<7)+(in_buffer[106]<<9))+(0-(in_buffer[107]<<0)-(in_buffer[107]<<2)-(in_buffer[107]<<4)+(in_buffer[107]<<8)+(in_buffer[107]<<9))-(0+(in_buffer[108]<<0)+(in_buffer[108]<<4)-(in_buffer[108]<<7)+(in_buffer[108]<<10))+(0+(in_buffer[109]<<0)-(in_buffer[109]<<3)+(in_buffer[109]<<8))+(0+(in_buffer[111]<<1)+(in_buffer[111]<<2)+(in_buffer[111]<<5)+(in_buffer[111]<<7))-(0+(in_buffer[112]<<1)-(in_buffer[112]<<4)+(in_buffer[112]<<9))+(0+(in_buffer[113]<<1)-(in_buffer[113]<<4)+(in_buffer[113]<<9))-(0+(in_buffer[114]<<0)-(in_buffer[114]<<3)+(in_buffer[114]<<8))+(0-(in_buffer[117]<<1)+(in_buffer[117]<<6)+(in_buffer[117]<<8)+(in_buffer[117]<<9))-(0+(in_buffer[118]<<2)+(in_buffer[118]<<3)+(in_buffer[118]<<6)+(in_buffer[118]<<8))+(0+(in_buffer[119]<<1)-(in_buffer[119]<<4)+(in_buffer[119]<<9))+(0+(in_buffer[120]<<0)+(in_buffer[120]<<2)+(in_buffer[120]<<6)+(in_buffer[120]<<9));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight17;
assign in_buffer_weight17=0-(0+(in_buffer[0]<<1)-(in_buffer[0]<<5)-(in_buffer[0]<<10)+(in_buffer[0]<<13))-(0-(in_buffer[1]<<0)-(in_buffer[1]<<3)+(in_buffer[1]<<6)+(in_buffer[1]<<10))-(0-(in_buffer[2]<<3)+(in_buffer[2]<<8)+(in_buffer[2]<<10)+(in_buffer[2]<<11))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<1)+(in_buffer[3]<<4)+(in_buffer[3]<<8)+(in_buffer[3]<<10)+(in_buffer[3]<<12))-(0+(in_buffer[4]<<4)+(in_buffer[4]<<5)+(in_buffer[4]<<8)+(in_buffer[4]<<10))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3)+(in_buffer[5]<<6)+(in_buffer[5]<<8)+(in_buffer[5]<<10)+(in_buffer[5]<<11))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<3)+(in_buffer[6]<<5)+(in_buffer[6]<<9)+(in_buffer[6]<<10))+(0+(in_buffer[7]<<2)-(in_buffer[7]<<4)-(in_buffer[7]<<7)+(in_buffer[7]<<10)+(in_buffer[7]<<12))+(0-(in_buffer[8]<<2)-(in_buffer[8]<<4)-(in_buffer[8]<<6)+(in_buffer[8]<<10)+(in_buffer[8]<<11))+(0-(in_buffer[9]<<1)-(in_buffer[9]<<3)-(in_buffer[9]<<5)+(in_buffer[9]<<9)+(in_buffer[9]<<10))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<3)+(in_buffer[10]<<5)+(in_buffer[10]<<9)+(in_buffer[10]<<10))+(0+(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<4)+(in_buffer[11]<<10)+(in_buffer[11]<<12))-(0+(in_buffer[12]<<1)-(in_buffer[12]<<3)-(in_buffer[12]<<6)+(in_buffer[12]<<9)+(in_buffer[12]<<11))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2)-(in_buffer[13]<<8)+(in_buffer[13]<<11)+(in_buffer[13]<<12))-(0-(in_buffer[14]<<1)-(in_buffer[14]<<4)+(in_buffer[14]<<7)+(in_buffer[14]<<11))+(0-(in_buffer[15]<<0)-(in_buffer[15]<<3)+(in_buffer[15]<<6)+(in_buffer[15]<<10))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<2)+(in_buffer[16]<<5)+(in_buffer[16]<<7))-(0+(in_buffer[17]<<2)-(in_buffer[17]<<5)+(in_buffer[17]<<10))+(0+(in_buffer[18]<<4)+(in_buffer[18]<<5)+(in_buffer[18]<<8)+(in_buffer[18]<<10))-(0-(in_buffer[19]<<0)+(in_buffer[19]<<4)-(in_buffer[19]<<6)-(in_buffer[19]<<8)+(in_buffer[19]<<11))+(0+(in_buffer[20]<<2)-(in_buffer[20]<<5)+(in_buffer[20]<<10))-(0+(in_buffer[21]<<3)+(in_buffer[21]<<4)+(in_buffer[21]<<7)+(in_buffer[21]<<9))+(0+(in_buffer[22]<<0)-(in_buffer[22]<<2)-(in_buffer[22]<<5)+(in_buffer[22]<<8)+(in_buffer[22]<<10))-(0+(in_buffer[23]<<2)-(in_buffer[23]<<5)+(in_buffer[23]<<10))+(0+(in_buffer[24]<<1)+(in_buffer[24]<<5)-(in_buffer[24]<<8)+(in_buffer[24]<<11))+(0-(in_buffer[25]<<0)-(in_buffer[25]<<2)-(in_buffer[25]<<4)+(in_buffer[25]<<8)+(in_buffer[25]<<9))-(0+(in_buffer[26]<<0)+(in_buffer[26]<<4)-(in_buffer[26]<<7)+(in_buffer[26]<<10))+(0+(in_buffer[27]<<0)+(in_buffer[27]<<2)+(in_buffer[27]<<4)-(in_buffer[27]<<6)+(in_buffer[27]<<9)+(in_buffer[27]<<12))-(0+(in_buffer[28]<<3)+(in_buffer[28]<<4)+(in_buffer[28]<<7)+(in_buffer[28]<<9))-(0-(in_buffer[29]<<0)+(in_buffer[29]<<10)+(in_buffer[29]<<11))-(0+(in_buffer[30]<<2)+(in_buffer[30]<<3)+(in_buffer[30]<<6)+(in_buffer[30]<<8))+(0-(in_buffer[31]<<0)-(in_buffer[31]<<3)+(in_buffer[31]<<6)+(in_buffer[31]<<10))-(0+(in_buffer[32]<<1)+(in_buffer[32]<<2)-(in_buffer[32]<<8)+(in_buffer[32]<<10)+(in_buffer[32]<<11))+(0+(in_buffer[33]<<2)+(in_buffer[33]<<3)+(in_buffer[33]<<6)+(in_buffer[33]<<8))+(0+(in_buffer[34]<<1)+(in_buffer[34]<<3)+(in_buffer[34]<<7)+(in_buffer[34]<<10))-(0+(in_buffer[35]<<1)-(in_buffer[35]<<4)+(in_buffer[35]<<9))+(0-(in_buffer[36]<<1)-(in_buffer[36]<<3)-(in_buffer[36]<<5)+(in_buffer[36]<<9)+(in_buffer[36]<<10))-(0-(in_buffer[37]<<2)+(in_buffer[37]<<7)+(in_buffer[37]<<9)+(in_buffer[37]<<10))+(0+(in_buffer[38]<<0)+(in_buffer[38]<<2)+(in_buffer[38]<<6)+(in_buffer[38]<<9))-(0+(in_buffer[39]<<2)+(in_buffer[39]<<6)-(in_buffer[39]<<9)+(in_buffer[39]<<12))-(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)-(in_buffer[40]<<4)+(in_buffer[40]<<8)+(in_buffer[40]<<9))-(0+(in_buffer[41]<<3)+(in_buffer[41]<<5)+(in_buffer[41]<<9)+(in_buffer[41]<<12))-(0+(in_buffer[42]<<2)+(in_buffer[42]<<3)+(in_buffer[42]<<6)+(in_buffer[42]<<8))+(0-(in_buffer[43]<<1)-(in_buffer[43]<<3)-(in_buffer[43]<<5)+(in_buffer[43]<<9)+(in_buffer[43]<<10))-(0+(in_buffer[44]<<0)-(in_buffer[44]<<2)-(in_buffer[44]<<5)+(in_buffer[44]<<8)+(in_buffer[44]<<10))-(0+(in_buffer[45]<<0)-(in_buffer[45]<<3)+(in_buffer[45]<<8))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<2)+(in_buffer[47]<<4)-(in_buffer[47]<<6)+(in_buffer[47]<<9)+(in_buffer[47]<<12))-(0-(in_buffer[48]<<1)+(in_buffer[48]<<4)-(in_buffer[48]<<6)+(in_buffer[48]<<8)+(in_buffer[48]<<9)+(in_buffer[48]<<12))-(0-(in_buffer[49]<<0)-(in_buffer[49]<<2)-(in_buffer[49]<<5)+(in_buffer[49]<<8)-(in_buffer[49]<<10)+(in_buffer[49]<<13))-(0+(in_buffer[50]<<1)+(in_buffer[50]<<3)+(in_buffer[50]<<7)+(in_buffer[50]<<10))+(0-(in_buffer[51]<<0)+(in_buffer[51]<<3)-(in_buffer[51]<<6)+(in_buffer[51]<<10)+(in_buffer[51]<<12))-(0+(in_buffer[52]<<0)+(in_buffer[52]<<2)-(in_buffer[52]<<8)+(in_buffer[52]<<11)+(in_buffer[52]<<12))+(0-(in_buffer[53]<<1)-(in_buffer[53]<<3)+(in_buffer[53]<<6)+(in_buffer[53]<<12))+(0+(in_buffer[54]<<1)+(in_buffer[54]<<4)+(in_buffer[54]<<8)+(in_buffer[54]<<13))+(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<5)+(in_buffer[55]<<11))-(0+(in_buffer[56]<<0)-(in_buffer[56]<<3)-(in_buffer[56]<<5)-(in_buffer[56]<<7)+(in_buffer[56]<<10)+(in_buffer[56]<<11))+(0+(in_buffer[57]<<0)-(in_buffer[57]<<3)-(in_buffer[57]<<5)-(in_buffer[57]<<7)+(in_buffer[57]<<10)+(in_buffer[57]<<11))+(0-(in_buffer[58]<<4)+(in_buffer[58]<<9)+(in_buffer[58]<<11)+(in_buffer[58]<<12))+(0+(in_buffer[59]<<0)+(in_buffer[59]<<2)+(in_buffer[59]<<3)+(in_buffer[59]<<9)+(in_buffer[59]<<11))-(0-(in_buffer[60]<<0)-(in_buffer[60]<<2)-(in_buffer[60]<<5)+(in_buffer[60]<<8)-(in_buffer[60]<<10)+(in_buffer[60]<<13))-(0+(in_buffer[61]<<1)+(in_buffer[61]<<2)-(in_buffer[61]<<8)+(in_buffer[61]<<10)+(in_buffer[61]<<11))+(0-(in_buffer[62]<<0)+(in_buffer[62]<<3)+(in_buffer[62]<<4)+(in_buffer[62]<<7)-(in_buffer[62]<<9)+(in_buffer[62]<<12))+(0+(in_buffer[63]<<0)+(in_buffer[63]<<1)+(in_buffer[63]<<4)+(in_buffer[63]<<6))+(0-(in_buffer[64]<<1)-(in_buffer[64]<<3)+(in_buffer[64]<<6)+(in_buffer[64]<<12))-(0-(in_buffer[65]<<1)+(in_buffer[65]<<6)+(in_buffer[65]<<8)+(in_buffer[65]<<9))+(0+(in_buffer[66]<<3)+(in_buffer[66]<<5)+(in_buffer[66]<<9)+(in_buffer[66]<<12))-(0-(in_buffer[67]<<1)+(in_buffer[67]<<3)+(in_buffer[67]<<4)+(in_buffer[67]<<7)+(in_buffer[67]<<9)+(in_buffer[67]<<11)+(in_buffer[67]<<12))+(0+(in_buffer[68]<<0)-(in_buffer[68]<<3)-(in_buffer[68]<<6)-(in_buffer[68]<<9)+(in_buffer[68]<<11)+(in_buffer[68]<<12))+(0-(in_buffer[69]<<1)-(in_buffer[69]<<3)+(in_buffer[69]<<6)+(in_buffer[69]<<12))+(0+(in_buffer[70]<<1)-(in_buffer[70]<<3)-(in_buffer[70]<<6)+(in_buffer[70]<<9)+(in_buffer[70]<<11))-(0+(in_buffer[71]<<1)+(in_buffer[71]<<2)-(in_buffer[71]<<6)+(in_buffer[71]<<13))+(0+(in_buffer[72]<<3)+(in_buffer[72]<<4)+(in_buffer[72]<<7)+(in_buffer[72]<<9))+(0-(in_buffer[73]<<1)-(in_buffer[73]<<3)+(in_buffer[73]<<6)+(in_buffer[73]<<12))-(0+(in_buffer[74]<<3)+(in_buffer[74]<<4)+(in_buffer[74]<<7)+(in_buffer[74]<<9))-(0+(in_buffer[75]<<0)+(in_buffer[75]<<1)-(in_buffer[75]<<7)+(in_buffer[75]<<9)+(in_buffer[75]<<10))-(0+(in_buffer[76]<<2)+(in_buffer[76]<<3)-(in_buffer[76]<<9)+(in_buffer[76]<<11)+(in_buffer[76]<<12))+(0+(in_buffer[77]<<0)-(in_buffer[77]<<7)-(in_buffer[77]<<9)+(in_buffer[77]<<13))-(0-(in_buffer[78]<<0)+(in_buffer[78]<<4)-(in_buffer[78]<<6)-(in_buffer[78]<<8)+(in_buffer[78]<<11))+(0+(in_buffer[79]<<1)+(in_buffer[79]<<4)+(in_buffer[79]<<6)+(in_buffer[79]<<10)+(in_buffer[79]<<11))+(0-(in_buffer[80]<<0)+(in_buffer[80]<<2)+(in_buffer[80]<<3)+(in_buffer[80]<<6)+(in_buffer[80]<<8)+(in_buffer[80]<<10)+(in_buffer[80]<<11))+(0-(in_buffer[81]<<1)+(in_buffer[81]<<4)-(in_buffer[81]<<6)+(in_buffer[81]<<8)+(in_buffer[81]<<9)+(in_buffer[81]<<12))-(0-(in_buffer[82]<<3)-(in_buffer[82]<<5)-(in_buffer[82]<<7)+(in_buffer[82]<<11)+(in_buffer[82]<<12))+(0+(in_buffer[83]<<5)+(in_buffer[83]<<6)+(in_buffer[83]<<9)+(in_buffer[83]<<11))+(0+(in_buffer[84]<<0)+(in_buffer[84]<<3)-(in_buffer[84]<<5)-(in_buffer[84]<<8)-(in_buffer[84]<<10)+(in_buffer[84]<<13))-(0+(in_buffer[85]<<1)+(in_buffer[85]<<2)-(in_buffer[85]<<8)+(in_buffer[85]<<10)+(in_buffer[85]<<11))-(0+(in_buffer[86]<<0)+(in_buffer[86]<<2)+(in_buffer[86]<<6)+(in_buffer[86]<<9))-(0-(in_buffer[87]<<0)+(in_buffer[87]<<4)-(in_buffer[87]<<6)-(in_buffer[87]<<8)+(in_buffer[87]<<11))-(0+(in_buffer[88]<<1)-(in_buffer[88]<<4)+(in_buffer[88]<<9))-(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)-(in_buffer[89]<<4)+(in_buffer[89]<<8)+(in_buffer[89]<<9))+(0-(in_buffer[90]<<1)-(in_buffer[90]<<3)+(in_buffer[90]<<6)+(in_buffer[90]<<12))+(0+(in_buffer[91]<<1)+(in_buffer[91]<<5)-(in_buffer[91]<<8)+(in_buffer[91]<<11))+(0+(in_buffer[92]<<1)+(in_buffer[92]<<5)-(in_buffer[92]<<8)+(in_buffer[92]<<11))-(0+(in_buffer[93]<<1)+(in_buffer[93]<<3)+(in_buffer[93]<<6)+(in_buffer[93]<<8)+(in_buffer[93]<<11)+(in_buffer[93]<<12))+(0-(in_buffer[94]<<1)-(in_buffer[94]<<3)+(in_buffer[94]<<6)+(in_buffer[94]<<12))+(0-(in_buffer[95]<<4)+(in_buffer[95]<<9)+(in_buffer[95]<<11)+(in_buffer[95]<<12))-(0+(in_buffer[96]<<3)+(in_buffer[96]<<4)+(in_buffer[96]<<7)+(in_buffer[96]<<9))+(0+(in_buffer[97]<<1)-(in_buffer[97]<<4)+(in_buffer[97]<<9))-(0+(in_buffer[98]<<2)-(in_buffer[98]<<4)-(in_buffer[98]<<7)+(in_buffer[98]<<10)+(in_buffer[98]<<12))-(0+(in_buffer[99]<<2)-(in_buffer[99]<<5)+(in_buffer[99]<<10))+(0-(in_buffer[100]<<2)+(in_buffer[100]<<7)+(in_buffer[100]<<9)+(in_buffer[100]<<10))-(0-(in_buffer[101]<<0)+(in_buffer[101]<<10)+(in_buffer[101]<<11))+(0-(in_buffer[102]<<0)+(in_buffer[102]<<5)+(in_buffer[102]<<7)+(in_buffer[102]<<8))+(0+(in_buffer[103]<<0)+(in_buffer[103]<<3)+(in_buffer[103]<<7)+(in_buffer[103]<<12))-(0+(in_buffer[104]<<0)+(in_buffer[104]<<2)+(in_buffer[104]<<4)-(in_buffer[104]<<6)+(in_buffer[104]<<9)+(in_buffer[104]<<12))+(0-(in_buffer[105]<<1)-(in_buffer[105]<<3)+(in_buffer[105]<<6)+(in_buffer[105]<<12))+(0+(in_buffer[106]<<1)+(in_buffer[106]<<3)-(in_buffer[106]<<5)-(in_buffer[106]<<8)+(in_buffer[106]<<12))-(0+(in_buffer[107]<<3)+(in_buffer[107]<<5)+(in_buffer[107]<<9)+(in_buffer[107]<<12))+(0+(in_buffer[108]<<3)-(in_buffer[108]<<6)+(in_buffer[108]<<11))-(0-(in_buffer[109]<<1)+(in_buffer[109]<<6)+(in_buffer[109]<<8)+(in_buffer[109]<<9))+(0+(in_buffer[110]<<2)+(in_buffer[110]<<3)+(in_buffer[110]<<6)+(in_buffer[110]<<8))+(0-(in_buffer[111]<<0)-(in_buffer[111]<<2)+(in_buffer[111]<<7)+(in_buffer[111]<<9)+(in_buffer[111]<<12))-(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)+(in_buffer[112]<<7)+(in_buffer[112]<<9)+(in_buffer[112]<<12))+(0+(in_buffer[113]<<1)-(in_buffer[113]<<3)-(in_buffer[113]<<5)+(in_buffer[113]<<8)+(in_buffer[113]<<11)+(in_buffer[113]<<13))+(0+(in_buffer[114]<<0)-(in_buffer[114]<<2)+(in_buffer[114]<<5)+(in_buffer[114]<<7)+(in_buffer[114]<<8)+(in_buffer[114]<<11)+(in_buffer[114]<<12))-(0+(in_buffer[115]<<1)-(in_buffer[115]<<4)-(in_buffer[115]<<7)-(in_buffer[115]<<10)+(in_buffer[115]<<12)+(in_buffer[115]<<13))+(0+(in_buffer[116]<<0)+(in_buffer[116]<<3)+(in_buffer[116]<<7)+(in_buffer[116]<<12))+(0-(in_buffer[117]<<0)-(in_buffer[117]<<2)-(in_buffer[117]<<5)+(in_buffer[117]<<8)-(in_buffer[117]<<10)+(in_buffer[117]<<13))-(0+(in_buffer[118]<<1)-(in_buffer[118]<<3)+(in_buffer[118]<<7)-(in_buffer[118]<<9)+(in_buffer[118]<<13))-(0+(in_buffer[119]<<4)+(in_buffer[119]<<5)+(in_buffer[119]<<8)+(in_buffer[119]<<10))+(0+(in_buffer[120]<<1)-(in_buffer[120]<<4)+(in_buffer[120]<<9));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight18;
assign in_buffer_weight18=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<1)+(in_buffer[0]<<4)+(in_buffer[0]<<7)-(in_buffer[0]<<9)+(in_buffer[0]<<14))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)-(in_buffer[1]<<6)-(in_buffer[1]<<10)+(in_buffer[1]<<12)+(in_buffer[1]<<13))+(0-(in_buffer[2]<<0)-(in_buffer[2]<<3)+(in_buffer[2]<<6)+(in_buffer[2]<<10))+(0-(in_buffer[3]<<1)+(in_buffer[3]<<5)+(in_buffer[3]<<6)+(in_buffer[3]<<9)+(in_buffer[3]<<13))-(0-(in_buffer[4]<<2)-(in_buffer[4]<<4)-(in_buffer[4]<<6)+(in_buffer[4]<<10)+(in_buffer[4]<<11))+(0+(in_buffer[5]<<1)+(in_buffer[5]<<2)-(in_buffer[5]<<8)+(in_buffer[5]<<10)+(in_buffer[5]<<11))-(0-(in_buffer[6]<<1)+(in_buffer[6]<<4)+(in_buffer[6]<<5)+(in_buffer[6]<<8)-(in_buffer[6]<<10)+(in_buffer[6]<<13))-(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)-(in_buffer[7]<<10)+(in_buffer[7]<<14))-(0+(in_buffer[8]<<0)+(in_buffer[8]<<1)+(in_buffer[8]<<4)+(in_buffer[8]<<6)+(in_buffer[8]<<8)+(in_buffer[8]<<9)+(in_buffer[8]<<12)+(in_buffer[8]<<14))-(0-(in_buffer[9]<<1)+(in_buffer[9]<<4)-(in_buffer[9]<<6)+(in_buffer[9]<<8)+(in_buffer[9]<<9)+(in_buffer[9]<<12))+(0+(in_buffer[10]<<4)+(in_buffer[10]<<5)+(in_buffer[10]<<8)+(in_buffer[10]<<10))-(0+(in_buffer[11]<<2)-(in_buffer[11]<<5)+(in_buffer[11]<<10))+(0-(in_buffer[12]<<0)+(in_buffer[12]<<3)-(in_buffer[12]<<6)+(in_buffer[12]<<10)+(in_buffer[12]<<12))+(0+(in_buffer[13]<<1)-(in_buffer[13]<<5)-(in_buffer[13]<<10)+(in_buffer[13]<<13))+(0+(in_buffer[14]<<0)-(in_buffer[14]<<3)+(in_buffer[14]<<7)+(in_buffer[14]<<9)+(in_buffer[14]<<11)+(in_buffer[14]<<13))+(0+(in_buffer[15]<<1)-(in_buffer[15]<<4)+(in_buffer[15]<<9))+(0+(in_buffer[16]<<0)-(in_buffer[16]<<2)+(in_buffer[16]<<10)+(in_buffer[16]<<13))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<6)+(in_buffer[17]<<7)+(in_buffer[17]<<11))+(0+(in_buffer[18]<<4)+(in_buffer[18]<<5)+(in_buffer[18]<<8)+(in_buffer[18]<<10))-(0+(in_buffer[19]<<0)+(in_buffer[19]<<2)-(in_buffer[19]<<8)+(in_buffer[19]<<11)+(in_buffer[19]<<12))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<1)-(in_buffer[20]<<6)+(in_buffer[20]<<10)+(in_buffer[20]<<14))-(0+(in_buffer[21]<<7)+(in_buffer[21]<<8)+(in_buffer[21]<<11)+(in_buffer[21]<<13))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<1)-(in_buffer[22]<<5)+(in_buffer[22]<<12))+(0+(in_buffer[23]<<6)+(in_buffer[23]<<7)+(in_buffer[23]<<10)+(in_buffer[23]<<12))+(0+(in_buffer[24]<<1)+(in_buffer[24]<<7)+(in_buffer[24]<<8)+(in_buffer[24]<<12))+(0-(in_buffer[25]<<0)-(in_buffer[25]<<2)+(in_buffer[25]<<7)+(in_buffer[25]<<9)+(in_buffer[25]<<12))+(0+(in_buffer[26]<<2)-(in_buffer[26]<<5)+(in_buffer[26]<<10))-(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)-(in_buffer[27]<<4)+(in_buffer[27]<<8)+(in_buffer[27]<<9))-(0+(in_buffer[28]<<1)+(in_buffer[28]<<2)-(in_buffer[28]<<8)+(in_buffer[28]<<10)+(in_buffer[28]<<11))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<2)-(in_buffer[29]<<4)-(in_buffer[29]<<7)+(in_buffer[29]<<11))-(0-(in_buffer[30]<<0)+(in_buffer[30]<<4)+(in_buffer[30]<<5)+(in_buffer[30]<<8)+(in_buffer[30]<<12))-(0+(in_buffer[31]<<1)+(in_buffer[31]<<3)+(in_buffer[31]<<6)+(in_buffer[31]<<8)+(in_buffer[31]<<11)+(in_buffer[31]<<12))-(0-(in_buffer[32]<<1)+(in_buffer[32]<<4)+(in_buffer[32]<<5)+(in_buffer[32]<<8)-(in_buffer[32]<<10)+(in_buffer[32]<<13))+(0+(in_buffer[33]<<5)+(in_buffer[33]<<6)+(in_buffer[33]<<9)+(in_buffer[33]<<11))+(0+(in_buffer[34]<<1)-(in_buffer[34]<<5)-(in_buffer[34]<<10)+(in_buffer[34]<<13))+(0-(in_buffer[35]<<4)+(in_buffer[35]<<9)+(in_buffer[35]<<11)+(in_buffer[35]<<12))+(0+(in_buffer[36]<<1)+(in_buffer[36]<<3)+(in_buffer[36]<<4)+(in_buffer[36]<<10)+(in_buffer[36]<<12))-(0-(in_buffer[37]<<1)+(in_buffer[37]<<5)-(in_buffer[37]<<7)-(in_buffer[37]<<9)+(in_buffer[37]<<12))-(0+(in_buffer[38]<<3)-(in_buffer[38]<<6)+(in_buffer[38]<<11))-(0+(in_buffer[39]<<0)+(in_buffer[39]<<1)-(in_buffer[39]<<5)+(in_buffer[39]<<12))-(0+(in_buffer[40]<<0)+(in_buffer[40]<<1)+(in_buffer[40]<<4)+(in_buffer[40]<<6))+(0-(in_buffer[41]<<0)+(in_buffer[41]<<2)+(in_buffer[41]<<3)+(in_buffer[41]<<6)+(in_buffer[41]<<8)+(in_buffer[41]<<10)+(in_buffer[41]<<11))-(0+(in_buffer[42]<<0)-(in_buffer[42]<<3)+(in_buffer[42]<<8))-(0+(in_buffer[43]<<0)+(in_buffer[43]<<1)-(in_buffer[43]<<4)-(in_buffer[43]<<6)-(in_buffer[43]<<8)+(in_buffer[43]<<10)+(in_buffer[43]<<11))+(0+(in_buffer[44]<<0)+(in_buffer[44]<<2)+(in_buffer[44]<<4)+(in_buffer[44]<<7)+(in_buffer[44]<<9)+(in_buffer[44]<<10)+(in_buffer[44]<<13))+(0-(in_buffer[45]<<4)+(in_buffer[45]<<9)+(in_buffer[45]<<11)+(in_buffer[45]<<12))+(0+(in_buffer[46]<<3)+(in_buffer[46]<<7)-(in_buffer[46]<<10)+(in_buffer[46]<<13))+(0+(in_buffer[47]<<1)+(in_buffer[47]<<3)+(in_buffer[47]<<5)-(in_buffer[47]<<7)+(in_buffer[47]<<10)+(in_buffer[47]<<13))+(0+(in_buffer[48]<<1)+(in_buffer[48]<<5)-(in_buffer[48]<<8)+(in_buffer[48]<<11))-(0+(in_buffer[49]<<2)+(in_buffer[49]<<3)+(in_buffer[49]<<6)+(in_buffer[49]<<8))-(0-(in_buffer[50]<<1)+(in_buffer[50]<<4)-(in_buffer[50]<<6)+(in_buffer[50]<<8)+(in_buffer[50]<<9)+(in_buffer[50]<<12))+(0+(in_buffer[51]<<1)+(in_buffer[51]<<3)+(in_buffer[51]<<7)+(in_buffer[51]<<10))+(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<5)+(in_buffer[52]<<11))-(0-(in_buffer[53]<<0)+(in_buffer[53]<<4)-(in_buffer[53]<<6)-(in_buffer[53]<<8)+(in_buffer[53]<<11))+(0+(in_buffer[54]<<3)+(in_buffer[54]<<4)+(in_buffer[54]<<7)+(in_buffer[54]<<9))-(0+(in_buffer[55]<<0)-(in_buffer[55]<<5)+(in_buffer[55]<<11)+(in_buffer[55]<<13))-(0+(in_buffer[56]<<0)-(in_buffer[56]<<2)+(in_buffer[56]<<6)-(in_buffer[56]<<8)+(in_buffer[56]<<12))+(0+(in_buffer[57]<<4)+(in_buffer[57]<<5)+(in_buffer[57]<<8)+(in_buffer[57]<<10))+(0-(in_buffer[58]<<0)+(in_buffer[58]<<6)+(in_buffer[58]<<7)+(in_buffer[58]<<13))-(0+(in_buffer[59]<<0)+(in_buffer[59]<<1)+(in_buffer[59]<<4)+(in_buffer[59]<<6))+(0-(in_buffer[60]<<1)-(in_buffer[60]<<3)-(in_buffer[60]<<5)+(in_buffer[60]<<9)+(in_buffer[60]<<10))-(0+(in_buffer[61]<<2)-(in_buffer[61]<<4)-(in_buffer[61]<<7)+(in_buffer[61]<<10)+(in_buffer[61]<<12))+(0+(in_buffer[62]<<0)+(in_buffer[62]<<3)+(in_buffer[62]<<5)+(in_buffer[62]<<9)+(in_buffer[62]<<10))-(0+(in_buffer[63]<<2)+(in_buffer[63]<<3)+(in_buffer[63]<<6)+(in_buffer[63]<<8))+(0+(in_buffer[65]<<5)+(in_buffer[65]<<6)+(in_buffer[65]<<9)+(in_buffer[65]<<11))-(0-(in_buffer[66]<<5)+(in_buffer[66]<<10)+(in_buffer[66]<<12)+(in_buffer[66]<<13))-(0+(in_buffer[67]<<0)+(in_buffer[67]<<2)+(in_buffer[67]<<3)-(in_buffer[67]<<6)-(in_buffer[67]<<8)+(in_buffer[67]<<13))-(0+(in_buffer[68]<<3)+(in_buffer[68]<<4)+(in_buffer[68]<<7)+(in_buffer[68]<<9))+(0+(in_buffer[69]<<1)+(in_buffer[69]<<2)-(in_buffer[69]<<6)+(in_buffer[69]<<13))+(0-(in_buffer[70]<<2)-(in_buffer[70]<<4)-(in_buffer[70]<<6)+(in_buffer[70]<<10)+(in_buffer[70]<<11))+(0-(in_buffer[71]<<0)+(in_buffer[71]<<4)+(in_buffer[71]<<5)+(in_buffer[71]<<8)+(in_buffer[71]<<12))-(0+(in_buffer[72]<<0)+(in_buffer[72]<<1)-(in_buffer[72]<<5)+(in_buffer[72]<<12))+(0+(in_buffer[73]<<1)+(in_buffer[73]<<5)-(in_buffer[73]<<8)+(in_buffer[73]<<11))-(0+(in_buffer[74]<<1)+(in_buffer[74]<<5)-(in_buffer[74]<<8)+(in_buffer[74]<<11))+(0+(in_buffer[75]<<0)+(in_buffer[75]<<1)-(in_buffer[75]<<4)-(in_buffer[75]<<6)-(in_buffer[75]<<8)+(in_buffer[75]<<10)+(in_buffer[75]<<11))-(0+(in_buffer[76]<<0)+(in_buffer[76]<<6)+(in_buffer[76]<<7)+(in_buffer[76]<<11))-(0-(in_buffer[77]<<1)-(in_buffer[77]<<3)+(in_buffer[77]<<6)+(in_buffer[77]<<12))-(0-(in_buffer[78]<<0)+(in_buffer[78]<<10)+(in_buffer[78]<<11))+(0-(in_buffer[79]<<1)-(in_buffer[79]<<3)+(in_buffer[79]<<6)+(in_buffer[79]<<12))+(0+(in_buffer[80]<<1)-(in_buffer[80]<<3)+(in_buffer[80]<<7)-(in_buffer[80]<<9)+(in_buffer[80]<<13))-(0-(in_buffer[81]<<0)+(in_buffer[81]<<5)+(in_buffer[81]<<7)+(in_buffer[81]<<8))+(0-(in_buffer[82]<<1)+(in_buffer[82]<<11)+(in_buffer[82]<<12))-(0-(in_buffer[83]<<0)+(in_buffer[83]<<10)+(in_buffer[83]<<11))+(0-(in_buffer[84]<<2)-(in_buffer[84]<<5)+(in_buffer[84]<<8)+(in_buffer[84]<<12))-(0+(in_buffer[86]<<1)+(in_buffer[86]<<2)+(in_buffer[86]<<5)+(in_buffer[86]<<7))+(0+(in_buffer[87]<<1)+(in_buffer[87]<<2)+(in_buffer[87]<<5)+(in_buffer[87]<<7))-(0+(in_buffer[88]<<0)+(in_buffer[88]<<2)-(in_buffer[88]<<4)-(in_buffer[88]<<7)+(in_buffer[88]<<11))+(0+(in_buffer[89]<<2)+(in_buffer[89]<<3)+(in_buffer[89]<<6)+(in_buffer[89]<<8))+(0+(in_buffer[90]<<1)+(in_buffer[90]<<3)+(in_buffer[90]<<4)+(in_buffer[90]<<10)+(in_buffer[90]<<12))+(0+(in_buffer[91]<<1)-(in_buffer[91]<<4)-(in_buffer[91]<<6)-(in_buffer[91]<<8)+(in_buffer[91]<<11)+(in_buffer[91]<<12))-(0-(in_buffer[92]<<0)-(in_buffer[92]<<3)+(in_buffer[92]<<8)+(in_buffer[92]<<11)+(in_buffer[92]<<12))+(0+(in_buffer[93]<<0)+(in_buffer[93]<<5)+(in_buffer[93]<<8)+(in_buffer[93]<<9)+(in_buffer[93]<<12))+(0+(in_buffer[94]<<1)+(in_buffer[94]<<3)-(in_buffer[94]<<5)-(in_buffer[94]<<8)+(in_buffer[94]<<12))+(0+(in_buffer[95]<<0)-(in_buffer[95]<<2)+(in_buffer[95]<<10)+(in_buffer[95]<<13))-(0+(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6)-(in_buffer[96]<<8)+(in_buffer[96]<<12))-(0+(in_buffer[97]<<1)+(in_buffer[97]<<3)+(in_buffer[97]<<6)+(in_buffer[97]<<8)+(in_buffer[97]<<11)+(in_buffer[97]<<12))-(0-(in_buffer[98]<<0)+(in_buffer[98]<<3)+(in_buffer[98]<<4)+(in_buffer[98]<<7)-(in_buffer[98]<<9)+(in_buffer[98]<<12))-(0-(in_buffer[99]<<0)+(in_buffer[99]<<4)-(in_buffer[99]<<6)-(in_buffer[99]<<8)+(in_buffer[99]<<11))-(0-(in_buffer[100]<<1)-(in_buffer[100]<<3)-(in_buffer[100]<<5)+(in_buffer[100]<<9)+(in_buffer[100]<<10))+(0+(in_buffer[101]<<0)-(in_buffer[101]<<2)+(in_buffer[101]<<6)-(in_buffer[101]<<8)+(in_buffer[101]<<12))+(0-(in_buffer[102]<<1)+(in_buffer[102]<<4)-(in_buffer[102]<<6)+(in_buffer[102]<<8)+(in_buffer[102]<<9)+(in_buffer[102]<<12))-(0+(in_buffer[103]<<0)-(in_buffer[103]<<2)+(in_buffer[103]<<6)-(in_buffer[103]<<8)+(in_buffer[103]<<12))+(0+(in_buffer[104]<<0)+(in_buffer[104]<<2)-(in_buffer[104]<<4)-(in_buffer[104]<<7)+(in_buffer[104]<<11))+(0-(in_buffer[105]<<3)+(in_buffer[105]<<8)+(in_buffer[105]<<10)+(in_buffer[105]<<11))+(0-(in_buffer[106]<<0)+(in_buffer[106]<<2)+(in_buffer[106]<<3)-(in_buffer[106]<<6)-(in_buffer[106]<<8)-(in_buffer[106]<<11)+(in_buffer[106]<<14))+(0+(in_buffer[107]<<0)+(in_buffer[107]<<3)+(in_buffer[107]<<5)+(in_buffer[107]<<9)+(in_buffer[107]<<10))-(0+(in_buffer[108]<<0)+(in_buffer[108]<<1)-(in_buffer[108]<<5)+(in_buffer[108]<<12))-(0+(in_buffer[109]<<0)+(in_buffer[109]<<1)-(in_buffer[109]<<4)-(in_buffer[109]<<6)-(in_buffer[109]<<8)+(in_buffer[109]<<10)+(in_buffer[109]<<11))+(0+(in_buffer[110]<<2)+(in_buffer[110]<<4)-(in_buffer[110]<<6)-(in_buffer[110]<<9)+(in_buffer[110]<<13))+(0+(in_buffer[111]<<0)+(in_buffer[111]<<1)-(in_buffer[111]<<7)+(in_buffer[111]<<9)+(in_buffer[111]<<10))-(0+(in_buffer[112]<<2)-(in_buffer[112]<<5)+(in_buffer[112]<<10))-(0+(in_buffer[113]<<0)+(in_buffer[113]<<2)+(in_buffer[113]<<3)-(in_buffer[113]<<6)-(in_buffer[113]<<8)+(in_buffer[113]<<13))-(0+(in_buffer[114]<<0)-(in_buffer[114]<<2)-(in_buffer[114]<<4)+(in_buffer[114]<<7)+(in_buffer[114]<<10)+(in_buffer[114]<<12))+(0+(in_buffer[115]<<1)+(in_buffer[115]<<2)-(in_buffer[115]<<6)+(in_buffer[115]<<13))+(0+(in_buffer[116]<<1)+(in_buffer[116]<<4)+(in_buffer[116]<<6)+(in_buffer[116]<<10)+(in_buffer[116]<<11))+(0+(in_buffer[117]<<2)+(in_buffer[117]<<8)+(in_buffer[117]<<9)+(in_buffer[117]<<13))+(0-(in_buffer[118]<<0)+(in_buffer[118]<<4)-(in_buffer[118]<<6)-(in_buffer[118]<<8)+(in_buffer[118]<<11))+(0+(in_buffer[119]<<0)+(in_buffer[119]<<4)+(in_buffer[119]<<6)+(in_buffer[119]<<11)+(in_buffer[119]<<12))+(0+(in_buffer[120]<<1)+(in_buffer[120]<<4)-(in_buffer[120]<<6)-(in_buffer[120]<<9)-(in_buffer[120]<<11)+(in_buffer[120]<<14));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight19;
assign in_buffer_weight19=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<3)-(in_buffer[0]<<6)+(in_buffer[0]<<10)+(in_buffer[0]<<12))-(0+(in_buffer[1]<<4)-(in_buffer[1]<<6)-(in_buffer[1]<<9)+(in_buffer[1]<<12)+(in_buffer[1]<<14))-(0+(in_buffer[2]<<2)+(in_buffer[2]<<4)+(in_buffer[2]<<6)-(in_buffer[2]<<8)+(in_buffer[2]<<11)+(in_buffer[2]<<14))-(0+(in_buffer[3]<<2)+(in_buffer[3]<<4)-(in_buffer[3]<<6)-(in_buffer[3]<<9)+(in_buffer[3]<<13))+(0-(in_buffer[4]<<1)-(in_buffer[4]<<3)-(in_buffer[4]<<5)+(in_buffer[4]<<9)+(in_buffer[4]<<10))+(0+(in_buffer[5]<<4)-(in_buffer[5]<<7)+(in_buffer[5]<<12))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<3)-(in_buffer[6]<<6)+(in_buffer[6]<<10)+(in_buffer[6]<<12))-(0-(in_buffer[7]<<2)-(in_buffer[7]<<5)+(in_buffer[7]<<8)+(in_buffer[7]<<12))-(0+(in_buffer[8]<<0)-(in_buffer[8]<<3)-(in_buffer[8]<<5)+(in_buffer[8]<<8)+(in_buffer[8]<<10)+(in_buffer[8]<<12)+(in_buffer[8]<<13))-(0-(in_buffer[9]<<1)-(in_buffer[9]<<3)+(in_buffer[9]<<8)+(in_buffer[9]<<10)+(in_buffer[9]<<13))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<4)-(in_buffer[10]<<7)+(in_buffer[10]<<10))-(0-(in_buffer[11]<<1)-(in_buffer[11]<<3)-(in_buffer[11]<<5)+(in_buffer[11]<<9)+(in_buffer[11]<<10))-(0+(in_buffer[12]<<3)+(in_buffer[12]<<4)+(in_buffer[12]<<7)+(in_buffer[12]<<9))-(0+(in_buffer[13]<<3)-(in_buffer[13]<<6)+(in_buffer[13]<<11))-(0-(in_buffer[14]<<1)-(in_buffer[14]<<3)+(in_buffer[14]<<6)+(in_buffer[14]<<12))-(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)+(in_buffer[15]<<5)+(in_buffer[15]<<11))+(0-(in_buffer[16]<<1)+(in_buffer[16]<<5)-(in_buffer[16]<<7)-(in_buffer[16]<<9)+(in_buffer[16]<<12))-(0-(in_buffer[17]<<0)-(in_buffer[17]<<3)+(in_buffer[17]<<6)+(in_buffer[17]<<10))-(0-(in_buffer[18]<<1)+(in_buffer[18]<<5)-(in_buffer[18]<<7)-(in_buffer[18]<<9)+(in_buffer[18]<<12))-(0+(in_buffer[19]<<5)+(in_buffer[19]<<6)+(in_buffer[19]<<9)+(in_buffer[19]<<11))+(0-(in_buffer[20]<<2)-(in_buffer[20]<<4)-(in_buffer[20]<<6)+(in_buffer[20]<<10)+(in_buffer[20]<<11))+(0+(in_buffer[21]<<1)-(in_buffer[21]<<5)-(in_buffer[21]<<10)+(in_buffer[21]<<13))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<4)+(in_buffer[22]<<6)+(in_buffer[22]<<11)+(in_buffer[22]<<12))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)-(in_buffer[23]<<8)+(in_buffer[23]<<11)+(in_buffer[23]<<12))+(0+(in_buffer[24]<<1)+(in_buffer[24]<<7)+(in_buffer[24]<<8)+(in_buffer[24]<<12))-(0-(in_buffer[25]<<0)+(in_buffer[25]<<4)-(in_buffer[25]<<6)-(in_buffer[25]<<8)+(in_buffer[25]<<11))-(0+(in_buffer[26]<<1)+(in_buffer[26]<<2)+(in_buffer[26]<<5)+(in_buffer[26]<<7))+(0-(in_buffer[27]<<1)-(in_buffer[27]<<3)-(in_buffer[27]<<5)+(in_buffer[27]<<9)+(in_buffer[27]<<10))+(0+(in_buffer[28]<<0)+(in_buffer[28]<<1)+(in_buffer[28]<<4)+(in_buffer[28]<<6))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)-(in_buffer[29]<<4)+(in_buffer[29]<<8)+(in_buffer[29]<<9))+(0+(in_buffer[30]<<0)+(in_buffer[30]<<1)-(in_buffer[30]<<5)+(in_buffer[30]<<12))+(0+(in_buffer[31]<<0)+(in_buffer[31]<<2)-(in_buffer[31]<<5)+(in_buffer[31]<<7)+(in_buffer[31]<<8)+(in_buffer[31]<<13))+(0-(in_buffer[32]<<1)+(in_buffer[32]<<5)+(in_buffer[32]<<6)+(in_buffer[32]<<9)+(in_buffer[32]<<13))-(0-(in_buffer[33]<<0)-(in_buffer[33]<<2)-(in_buffer[33]<<4)-(in_buffer[33]<<6)+(in_buffer[33]<<11)+(in_buffer[33]<<12))+(0+(in_buffer[34]<<4)+(in_buffer[34]<<5)+(in_buffer[34]<<8)+(in_buffer[34]<<10))+(0+(in_buffer[35]<<5)+(in_buffer[35]<<6)+(in_buffer[35]<<9)+(in_buffer[35]<<11))-(0-(in_buffer[36]<<2)-(in_buffer[36]<<4)-(in_buffer[36]<<6)+(in_buffer[36]<<10)+(in_buffer[36]<<11))-(0+(in_buffer[37]<<1)+(in_buffer[37]<<2)+(in_buffer[37]<<5)+(in_buffer[37]<<7))-(0+(in_buffer[38]<<0)-(in_buffer[38]<<4)-(in_buffer[38]<<9)+(in_buffer[38]<<12))+(0+(in_buffer[39]<<1)-(in_buffer[39]<<4)+(in_buffer[39]<<9))+(0+(in_buffer[42]<<1)-(in_buffer[42]<<5)-(in_buffer[42]<<10)+(in_buffer[42]<<13))-(0+(in_buffer[43]<<0)+(in_buffer[43]<<1)+(in_buffer[43]<<4)+(in_buffer[43]<<6))-(0+(in_buffer[44]<<0)+(in_buffer[44]<<2)-(in_buffer[44]<<6)-(in_buffer[44]<<10)+(in_buffer[44]<<12)+(in_buffer[44]<<13))-(0-(in_buffer[45]<<1)-(in_buffer[45]<<4)+(in_buffer[45]<<7)+(in_buffer[45]<<11))+(0-(in_buffer[46]<<0)+(in_buffer[46]<<2)+(in_buffer[46]<<3)+(in_buffer[46]<<6)+(in_buffer[46]<<8)+(in_buffer[46]<<10)+(in_buffer[46]<<11))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<1)-(in_buffer[47]<<7)+(in_buffer[47]<<9)+(in_buffer[47]<<10))+(0-(in_buffer[48]<<0)-(in_buffer[48]<<2)-(in_buffer[48]<<4)+(in_buffer[48]<<8)+(in_buffer[48]<<9))-(0+(in_buffer[49]<<0)+(in_buffer[49]<<4)-(in_buffer[49]<<7)+(in_buffer[49]<<10))+(0+(in_buffer[50]<<0)+(in_buffer[50]<<6)+(in_buffer[50]<<7)+(in_buffer[50]<<11))+(0-(in_buffer[51]<<0)-(in_buffer[51]<<2)+(in_buffer[51]<<7)+(in_buffer[51]<<9)+(in_buffer[51]<<12))+(0-(in_buffer[52]<<0)+(in_buffer[52]<<4)-(in_buffer[52]<<6)-(in_buffer[52]<<8)+(in_buffer[52]<<11))+(0-(in_buffer[53]<<0)+(in_buffer[53]<<3)-(in_buffer[53]<<5)+(in_buffer[53]<<7)+(in_buffer[53]<<8)+(in_buffer[53]<<11))-(0+(in_buffer[54]<<4)-(in_buffer[54]<<7)+(in_buffer[54]<<12))-(0+(in_buffer[55]<<0)-(in_buffer[55]<<5)+(in_buffer[55]<<11)+(in_buffer[55]<<13))+(0-(in_buffer[56]<<0)-(in_buffer[56]<<2)+(in_buffer[56]<<7)+(in_buffer[56]<<9)+(in_buffer[56]<<12))+(0+(in_buffer[57]<<1)-(in_buffer[57]<<4)+(in_buffer[57]<<9))+(0+(in_buffer[58]<<2)-(in_buffer[58]<<5)+(in_buffer[58]<<10))+(0-(in_buffer[59]<<0)-(in_buffer[59]<<3)+(in_buffer[59]<<6)+(in_buffer[59]<<10))+(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)+(in_buffer[60]<<4)+(in_buffer[60]<<6))+(0-(in_buffer[61]<<0)-(in_buffer[61]<<2)-(in_buffer[61]<<4)+(in_buffer[61]<<8)+(in_buffer[61]<<9))+(0+(in_buffer[62]<<1)-(in_buffer[62]<<3)-(in_buffer[62]<<6)+(in_buffer[62]<<9)+(in_buffer[62]<<11))+(0-(in_buffer[63]<<1)+(in_buffer[63]<<6)+(in_buffer[63]<<8)+(in_buffer[63]<<9))-(0-(in_buffer[64]<<0)+(in_buffer[64]<<5)+(in_buffer[64]<<7)+(in_buffer[64]<<8))-(0+(in_buffer[65]<<1)-(in_buffer[65]<<4)-(in_buffer[65]<<6)-(in_buffer[65]<<8)+(in_buffer[65]<<11)+(in_buffer[65]<<12))-(0-(in_buffer[66]<<1)+(in_buffer[66]<<6)+(in_buffer[66]<<8)+(in_buffer[66]<<9))+(0-(in_buffer[67]<<0)+(in_buffer[67]<<4)+(in_buffer[67]<<5)+(in_buffer[67]<<8)+(in_buffer[67]<<12))-(0+(in_buffer[68]<<0)+(in_buffer[68]<<1)+(in_buffer[68]<<4)+(in_buffer[68]<<6))+(0+(in_buffer[69]<<0)+(in_buffer[69]<<1)-(in_buffer[69]<<7)+(in_buffer[69]<<9)+(in_buffer[69]<<10))-(0+(in_buffer[71]<<2)-(in_buffer[71]<<5)+(in_buffer[71]<<10))+(0+(in_buffer[72]<<3)+(in_buffer[72]<<4)+(in_buffer[72]<<7)+(in_buffer[72]<<9))+(0-(in_buffer[73]<<0)-(in_buffer[73]<<2)-(in_buffer[73]<<4)+(in_buffer[73]<<8)+(in_buffer[73]<<9))+(0+(in_buffer[74]<<3)+(in_buffer[74]<<4)+(in_buffer[74]<<7)+(in_buffer[74]<<9))-(0+(in_buffer[75]<<0)-(in_buffer[75]<<3)+(in_buffer[75]<<8))-(0-(in_buffer[76]<<0)+(in_buffer[76]<<2)+(in_buffer[76]<<3)+(in_buffer[76]<<6)+(in_buffer[76]<<8)+(in_buffer[76]<<10)+(in_buffer[76]<<11))+(0+(in_buffer[77]<<1)+(in_buffer[77]<<3)+(in_buffer[77]<<7)+(in_buffer[77]<<10))+(0-(in_buffer[78]<<0)-(in_buffer[78]<<3)+(in_buffer[78]<<6)+(in_buffer[78]<<10))-(0+(in_buffer[79]<<0)-(in_buffer[79]<<3)-(in_buffer[79]<<5)-(in_buffer[79]<<7)+(in_buffer[79]<<10)+(in_buffer[79]<<11))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<3)+(in_buffer[80]<<6)+(in_buffer[80]<<10))+(0+(in_buffer[81]<<0)+(in_buffer[81]<<6)+(in_buffer[81]<<7)+(in_buffer[81]<<11))+(0+(in_buffer[82]<<0)-(in_buffer[82]<<3)-(in_buffer[82]<<5)-(in_buffer[82]<<7)+(in_buffer[82]<<10)+(in_buffer[82]<<11))+(0+(in_buffer[83]<<0)-(in_buffer[83]<<3)+(in_buffer[83]<<8))+(0+(in_buffer[84]<<2)+(in_buffer[84]<<3)+(in_buffer[84]<<6)+(in_buffer[84]<<8))-(0+(in_buffer[85]<<0)-(in_buffer[85]<<2)-(in_buffer[85]<<5)+(in_buffer[85]<<8)+(in_buffer[85]<<10))-(0+(in_buffer[86]<<4)+(in_buffer[86]<<5)+(in_buffer[86]<<8)+(in_buffer[86]<<10))-(0-(in_buffer[87]<<2)-(in_buffer[87]<<5)+(in_buffer[87]<<8)+(in_buffer[87]<<12))+(0-(in_buffer[88]<<0)+(in_buffer[88]<<4)-(in_buffer[88]<<6)-(in_buffer[88]<<8)+(in_buffer[88]<<11))+(0+(in_buffer[89]<<0)+(in_buffer[89]<<2)+(in_buffer[89]<<3)+(in_buffer[89]<<9)+(in_buffer[89]<<11))-(0-(in_buffer[90]<<1)-(in_buffer[90]<<3)+(in_buffer[90]<<6)+(in_buffer[90]<<12))-(0-(in_buffer[91]<<0)+(in_buffer[91]<<3)+(in_buffer[91]<<4)+(in_buffer[91]<<7)-(in_buffer[91]<<9)+(in_buffer[91]<<12))+(0+(in_buffer[92]<<1)+(in_buffer[92]<<5)-(in_buffer[92]<<8)+(in_buffer[92]<<11))+(0-(in_buffer[93]<<0)+(in_buffer[93]<<4)-(in_buffer[93]<<6)-(in_buffer[93]<<8)+(in_buffer[93]<<11))-(0+(in_buffer[94]<<0)+(in_buffer[94]<<1)-(in_buffer[94]<<7)+(in_buffer[94]<<9)+(in_buffer[94]<<10))-(0+(in_buffer[95]<<0)+(in_buffer[95]<<5)+(in_buffer[95]<<8)+(in_buffer[95]<<9)+(in_buffer[95]<<12))-(0+(in_buffer[96]<<0)-(in_buffer[96]<<2)+(in_buffer[96]<<6)-(in_buffer[96]<<8)+(in_buffer[96]<<12))-(0-(in_buffer[97]<<1)+(in_buffer[97]<<6)+(in_buffer[97]<<8)+(in_buffer[97]<<9))-(0+(in_buffer[98]<<0)+(in_buffer[98]<<2)+(in_buffer[98]<<4)-(in_buffer[98]<<6)+(in_buffer[98]<<9)+(in_buffer[98]<<12))-(0+(in_buffer[99]<<5)-(in_buffer[99]<<8)+(in_buffer[99]<<13))+(0+(in_buffer[100]<<0)+(in_buffer[100]<<5)+(in_buffer[100]<<8)+(in_buffer[100]<<9)+(in_buffer[100]<<12))-(0+(in_buffer[101]<<2)+(in_buffer[101]<<4)+(in_buffer[101]<<8)+(in_buffer[101]<<11))-(0-(in_buffer[102]<<0)+(in_buffer[102]<<3)-(in_buffer[102]<<5)+(in_buffer[102]<<7)+(in_buffer[102]<<8)+(in_buffer[102]<<11))+(0+(in_buffer[103]<<3)-(in_buffer[103]<<6)+(in_buffer[103]<<11))-(0+(in_buffer[104]<<1)+(in_buffer[104]<<3)+(in_buffer[104]<<7)+(in_buffer[104]<<10))-(0-(in_buffer[105]<<0)-(in_buffer[105]<<3)+(in_buffer[105]<<6)+(in_buffer[105]<<10))-(0-(in_buffer[106]<<0)-(in_buffer[106]<<2)+(in_buffer[106]<<7)+(in_buffer[106]<<9)+(in_buffer[106]<<12))-(0-(in_buffer[107]<<2)-(in_buffer[107]<<4)-(in_buffer[107]<<6)+(in_buffer[107]<<10)+(in_buffer[107]<<11))-(0+(in_buffer[108]<<0)+(in_buffer[108]<<4)-(in_buffer[108]<<7)+(in_buffer[108]<<10))-(0-(in_buffer[109]<<1)+(in_buffer[109]<<4)-(in_buffer[109]<<7)+(in_buffer[109]<<11)+(in_buffer[109]<<13))-(0+(in_buffer[110]<<2)-(in_buffer[110]<<4)+(in_buffer[110]<<8)-(in_buffer[110]<<10)+(in_buffer[110]<<14))+(0-(in_buffer[111]<<2)+(in_buffer[111]<<6)-(in_buffer[111]<<8)-(in_buffer[111]<<10)+(in_buffer[111]<<13))+(0+(in_buffer[112]<<1)+(in_buffer[112]<<3)+(in_buffer[112]<<6)+(in_buffer[112]<<8)+(in_buffer[112]<<11)+(in_buffer[112]<<12))+(0+(in_buffer[113]<<2)+(in_buffer[113]<<3)+(in_buffer[113]<<6)+(in_buffer[113]<<8))-(0-(in_buffer[114]<<2)+(in_buffer[114]<<12)+(in_buffer[114]<<13))-(0+(in_buffer[115]<<1)+(in_buffer[115]<<2)-(in_buffer[115]<<5)-(in_buffer[115]<<8)+(in_buffer[115]<<14))-(0-(in_buffer[116]<<1)-(in_buffer[116]<<3)-(in_buffer[116]<<5)-(in_buffer[116]<<7)+(in_buffer[116]<<12)+(in_buffer[116]<<13))-(0-(in_buffer[117]<<0)-(in_buffer[117]<<2)+(in_buffer[117]<<7)+(in_buffer[117]<<9)+(in_buffer[117]<<12))+(0-(in_buffer[118]<<1)+(in_buffer[118]<<3)+(in_buffer[118]<<4)+(in_buffer[118]<<7)+(in_buffer[118]<<9)+(in_buffer[118]<<11)+(in_buffer[118]<<12))+(0-(in_buffer[119]<<2)-(in_buffer[119]<<5)+(in_buffer[119]<<8)+(in_buffer[119]<<12))-(0+(in_buffer[120]<<0)+(in_buffer[120]<<6)+(in_buffer[120]<<9)+(in_buffer[120]<<12)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight20;
assign in_buffer_weight20=0-(0+(in_buffer[0]<<5)-(in_buffer[0]<<8)+(in_buffer[0]<<13))-(0-(in_buffer[1]<<0)+(in_buffer[1]<<3)+(in_buffer[1]<<4)+(in_buffer[1]<<7)-(in_buffer[1]<<9)+(in_buffer[1]<<12))-(0+(in_buffer[2]<<0)-(in_buffer[2]<<2)-(in_buffer[2]<<4)+(in_buffer[2]<<7)+(in_buffer[2]<<10)+(in_buffer[2]<<12))+(0-(in_buffer[3]<<2)+(in_buffer[3]<<7)+(in_buffer[3]<<9)+(in_buffer[3]<<10))+(0+(in_buffer[4]<<5)+(in_buffer[4]<<6)+(in_buffer[4]<<9)+(in_buffer[4]<<11))+(0-(in_buffer[5]<<0)+(in_buffer[5]<<5)+(in_buffer[5]<<7)+(in_buffer[5]<<8))+(0+(in_buffer[6]<<4)-(in_buffer[6]<<7)+(in_buffer[6]<<12))+(0+(in_buffer[7]<<0)-(in_buffer[7]<<4)-(in_buffer[7]<<9)+(in_buffer[7]<<12))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<5)+(in_buffer[8]<<7)+(in_buffer[8]<<8))+(0-(in_buffer[9]<<1)-(in_buffer[9]<<4)+(in_buffer[9]<<7)+(in_buffer[9]<<11))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)-(in_buffer[10]<<4)-(in_buffer[10]<<6)-(in_buffer[10]<<8)+(in_buffer[10]<<10)+(in_buffer[10]<<11))-(0+(in_buffer[11]<<2)+(in_buffer[11]<<4)+(in_buffer[11]<<5)+(in_buffer[11]<<11)+(in_buffer[11]<<13))+(0-(in_buffer[12]<<1)+(in_buffer[12]<<4)+(in_buffer[12]<<5)+(in_buffer[12]<<8)-(in_buffer[12]<<10)+(in_buffer[12]<<13))+(0+(in_buffer[13]<<1)+(in_buffer[13]<<3)+(in_buffer[13]<<6)+(in_buffer[13]<<8)+(in_buffer[13]<<11)+(in_buffer[13]<<12))+(0-(in_buffer[14]<<0)+(in_buffer[14]<<5)+(in_buffer[14]<<7)+(in_buffer[14]<<8))-(0-(in_buffer[15]<<0)-(in_buffer[15]<<2)-(in_buffer[15]<<4)+(in_buffer[15]<<8)+(in_buffer[15]<<9))-(0-(in_buffer[16]<<0)-(in_buffer[16]<<2)-(in_buffer[16]<<4)-(in_buffer[16]<<6)+(in_buffer[16]<<11)+(in_buffer[16]<<12))-(0+(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<8)+(in_buffer[17]<<11))-(0+(in_buffer[18]<<0)+(in_buffer[18]<<3)+(in_buffer[18]<<7)+(in_buffer[18]<<12))+(0+(in_buffer[19]<<0)-(in_buffer[19]<<2)-(in_buffer[19]<<5)+(in_buffer[19]<<8)+(in_buffer[19]<<10))+(0+(in_buffer[20]<<5)-(in_buffer[20]<<8)+(in_buffer[20]<<13))-(0+(in_buffer[21]<<1)+(in_buffer[21]<<5)-(in_buffer[21]<<8)+(in_buffer[21]<<11))-(0-(in_buffer[22]<<0)+(in_buffer[22]<<4)+(in_buffer[22]<<6)+(in_buffer[22]<<12)+(in_buffer[22]<<13))+(0-(in_buffer[23]<<2)-(in_buffer[23]<<5)+(in_buffer[23]<<8)+(in_buffer[23]<<12))+(0-(in_buffer[24]<<1)+(in_buffer[24]<<5)-(in_buffer[24]<<7)-(in_buffer[24]<<9)+(in_buffer[24]<<12))+(0+(in_buffer[25]<<1)+(in_buffer[25]<<3)+(in_buffer[25]<<7)+(in_buffer[25]<<10))+(0+(in_buffer[26]<<0)+(in_buffer[26]<<1)+(in_buffer[26]<<4)+(in_buffer[26]<<6))-(0-(in_buffer[27]<<0)+(in_buffer[27]<<4)-(in_buffer[27]<<7)-(in_buffer[27]<<10)+(in_buffer[27]<<13))+(0-(in_buffer[28]<<0)+(in_buffer[28]<<5)+(in_buffer[28]<<7)+(in_buffer[28]<<8))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<3)+(in_buffer[29]<<6)+(in_buffer[29]<<10))+(0-(in_buffer[30]<<1)+(in_buffer[30]<<6)+(in_buffer[30]<<8)+(in_buffer[30]<<9))+(0+(in_buffer[31]<<2)+(in_buffer[31]<<4)+(in_buffer[31]<<8)+(in_buffer[31]<<11))-(0+(in_buffer[32]<<2)+(in_buffer[32]<<3)+(in_buffer[32]<<6)+(in_buffer[32]<<8))-(0-(in_buffer[33]<<1)-(in_buffer[33]<<3)+(in_buffer[33]<<6)+(in_buffer[33]<<12))+(0+(in_buffer[34]<<3)-(in_buffer[34]<<6)+(in_buffer[34]<<11))+(0-(in_buffer[35]<<1)-(in_buffer[35]<<4)+(in_buffer[35]<<7)+(in_buffer[35]<<11))-(0+(in_buffer[36]<<0)+(in_buffer[36]<<1)+(in_buffer[36]<<6)+(in_buffer[36]<<9)+(in_buffer[36]<<11)+(in_buffer[36]<<12))+(0-(in_buffer[37]<<2)-(in_buffer[37]<<4)-(in_buffer[37]<<6)+(in_buffer[37]<<10)+(in_buffer[37]<<11))-(0+(in_buffer[38]<<2)+(in_buffer[38]<<3)+(in_buffer[38]<<6)+(in_buffer[38]<<8))+(0-(in_buffer[39]<<1)-(in_buffer[39]<<3)+(in_buffer[39]<<6)+(in_buffer[39]<<12))-(0-(in_buffer[40]<<1)-(in_buffer[40]<<3)-(in_buffer[40]<<5)+(in_buffer[40]<<9)+(in_buffer[40]<<10))+(0-(in_buffer[41]<<1)-(in_buffer[41]<<3)+(in_buffer[41]<<6)+(in_buffer[41]<<12))-(0-(in_buffer[42]<<0)+(in_buffer[42]<<3)-(in_buffer[42]<<5)+(in_buffer[42]<<7)+(in_buffer[42]<<8)+(in_buffer[42]<<11))+(0-(in_buffer[43]<<1)+(in_buffer[43]<<3)+(in_buffer[43]<<4)+(in_buffer[43]<<7)+(in_buffer[43]<<9)+(in_buffer[43]<<11)+(in_buffer[43]<<12))-(0+(in_buffer[44]<<0)+(in_buffer[44]<<1)-(in_buffer[44]<<5)+(in_buffer[44]<<12))-(0+(in_buffer[45]<<0)+(in_buffer[45]<<2)+(in_buffer[45]<<6)+(in_buffer[45]<<9))+(0+(in_buffer[46]<<0)+(in_buffer[46]<<2)+(in_buffer[46]<<6)+(in_buffer[46]<<9))-(0+(in_buffer[47]<<0)-(in_buffer[47]<<7)-(in_buffer[47]<<9)+(in_buffer[47]<<13))+(0+(in_buffer[48]<<0)-(in_buffer[48]<<2)+(in_buffer[48]<<5)+(in_buffer[48]<<7)+(in_buffer[48]<<8)+(in_buffer[48]<<11)+(in_buffer[48]<<12))-(0-(in_buffer[49]<<0)+(in_buffer[49]<<5)+(in_buffer[49]<<7)+(in_buffer[49]<<8))-(0+(in_buffer[51]<<2)+(in_buffer[51]<<5)+(in_buffer[51]<<7)+(in_buffer[51]<<11)+(in_buffer[51]<<12))-(0+(in_buffer[52]<<1)-(in_buffer[52]<<4)+(in_buffer[52]<<9))-(0+(in_buffer[53]<<0)+(in_buffer[53]<<2)+(in_buffer[53]<<3)-(in_buffer[53]<<6)-(in_buffer[53]<<8)+(in_buffer[53]<<13))+(0+(in_buffer[54]<<1)+(in_buffer[54]<<7)+(in_buffer[54]<<8)+(in_buffer[54]<<12))-(0+(in_buffer[55]<<7)+(in_buffer[55]<<8)+(in_buffer[55]<<11)+(in_buffer[55]<<13))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<1)-(in_buffer[56]<<4)-(in_buffer[56]<<6)-(in_buffer[56]<<8)+(in_buffer[56]<<10)+(in_buffer[56]<<11))-(0+(in_buffer[57]<<0)-(in_buffer[57]<<3)+(in_buffer[57]<<8))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<1)-(in_buffer[58]<<5)+(in_buffer[58]<<12))+(0-(in_buffer[59]<<0)+(in_buffer[59]<<10)+(in_buffer[59]<<11))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)-(in_buffer[60]<<7)+(in_buffer[60]<<9)+(in_buffer[60]<<10))-(0+(in_buffer[61]<<2)+(in_buffer[61]<<4)+(in_buffer[61]<<8)+(in_buffer[61]<<11))-(0-(in_buffer[62]<<1)+(in_buffer[62]<<3)+(in_buffer[62]<<4)+(in_buffer[62]<<7)+(in_buffer[62]<<9)+(in_buffer[62]<<11)+(in_buffer[62]<<12))-(0+(in_buffer[63]<<0)+(in_buffer[63]<<2)-(in_buffer[63]<<4)-(in_buffer[63]<<7)+(in_buffer[63]<<11))+(0+(in_buffer[64]<<1)+(in_buffer[64]<<3)+(in_buffer[64]<<7)+(in_buffer[64]<<10))+(0+(in_buffer[65]<<0)+(in_buffer[65]<<6)+(in_buffer[65]<<9)+(in_buffer[65]<<12)+(in_buffer[65]<<13))-(0+(in_buffer[66]<<2)+(in_buffer[66]<<4)+(in_buffer[66]<<6)-(in_buffer[66]<<8)+(in_buffer[66]<<11)+(in_buffer[66]<<14))-(0+(in_buffer[67]<<0)+(in_buffer[67]<<2)+(in_buffer[67]<<4)-(in_buffer[67]<<6)+(in_buffer[67]<<9)+(in_buffer[67]<<12))+(0+(in_buffer[68]<<1)+(in_buffer[68]<<5)-(in_buffer[68]<<8)+(in_buffer[68]<<11))-(0+(in_buffer[69]<<0)-(in_buffer[69]<<2)-(in_buffer[69]<<5)+(in_buffer[69]<<8)+(in_buffer[69]<<10))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<4)-(in_buffer[70]<<7)+(in_buffer[70]<<10))+(0+(in_buffer[71]<<0)+(in_buffer[71]<<2)+(in_buffer[71]<<6)+(in_buffer[71]<<9))+(0-(in_buffer[72]<<1)+(in_buffer[72]<<6)+(in_buffer[72]<<8)+(in_buffer[72]<<9))-(0+(in_buffer[73]<<4)-(in_buffer[73]<<7)+(in_buffer[73]<<12))-(0-(in_buffer[74]<<0)-(in_buffer[74]<<3)+(in_buffer[74]<<6)+(in_buffer[74]<<10))+(0+(in_buffer[75]<<1)+(in_buffer[75]<<3)+(in_buffer[75]<<7)+(in_buffer[75]<<10))+(0-(in_buffer[76]<<1)+(in_buffer[76]<<5)-(in_buffer[76]<<7)-(in_buffer[76]<<9)+(in_buffer[76]<<12))-(0+(in_buffer[77]<<2)-(in_buffer[77]<<4)-(in_buffer[77]<<7)+(in_buffer[77]<<10)+(in_buffer[77]<<12))-(0+(in_buffer[78]<<0)+(in_buffer[78]<<2)+(in_buffer[78]<<4)-(in_buffer[78]<<6)+(in_buffer[78]<<9)+(in_buffer[78]<<12))+(0+(in_buffer[79]<<1)+(in_buffer[79]<<2)-(in_buffer[79]<<5)-(in_buffer[79]<<7)-(in_buffer[79]<<9)+(in_buffer[79]<<11)+(in_buffer[79]<<12))+(0+(in_buffer[80]<<3)+(in_buffer[80]<<4)+(in_buffer[80]<<7)+(in_buffer[80]<<9))+(0+(in_buffer[81]<<0)+(in_buffer[81]<<1)-(in_buffer[81]<<4)-(in_buffer[81]<<6)-(in_buffer[81]<<8)+(in_buffer[81]<<10)+(in_buffer[81]<<11))+(0+(in_buffer[82]<<0)-(in_buffer[82]<<3)-(in_buffer[82]<<5)-(in_buffer[82]<<7)+(in_buffer[82]<<10)+(in_buffer[82]<<11))+(0-(in_buffer[83]<<1)+(in_buffer[83]<<5)-(in_buffer[83]<<7)-(in_buffer[83]<<9)+(in_buffer[83]<<12))-(0+(in_buffer[84]<<0)+(in_buffer[84]<<2)-(in_buffer[84]<<4)-(in_buffer[84]<<7)+(in_buffer[84]<<11))+(0+(in_buffer[85]<<0)-(in_buffer[85]<<2)-(in_buffer[85]<<5)+(in_buffer[85]<<8)+(in_buffer[85]<<10))+(0-(in_buffer[86]<<2)+(in_buffer[86]<<7)+(in_buffer[86]<<9)+(in_buffer[86]<<10))-(0+(in_buffer[87]<<1)+(in_buffer[87]<<2)-(in_buffer[87]<<5)-(in_buffer[87]<<7)-(in_buffer[87]<<9)+(in_buffer[87]<<11)+(in_buffer[87]<<12))-(0-(in_buffer[88]<<0)+(in_buffer[88]<<4)-(in_buffer[88]<<7)-(in_buffer[88]<<10)+(in_buffer[88]<<13))-(0-(in_buffer[89]<<0)-(in_buffer[89]<<3)+(in_buffer[89]<<6)+(in_buffer[89]<<10))-(0+(in_buffer[90]<<0)-(in_buffer[90]<<2)-(in_buffer[90]<<5)+(in_buffer[90]<<8)+(in_buffer[90]<<10))-(0-(in_buffer[91]<<0)-(in_buffer[91]<<2)-(in_buffer[91]<<4)+(in_buffer[91]<<8)+(in_buffer[91]<<9))+(0-(in_buffer[92]<<0)+(in_buffer[92]<<2)+(in_buffer[92]<<3)+(in_buffer[92]<<6)+(in_buffer[92]<<8)+(in_buffer[92]<<10)+(in_buffer[92]<<11))+(0-(in_buffer[93]<<0)+(in_buffer[93]<<2)+(in_buffer[93]<<3)+(in_buffer[93]<<6)+(in_buffer[93]<<8)+(in_buffer[93]<<10)+(in_buffer[93]<<11))+(0+(in_buffer[94]<<0)+(in_buffer[94]<<2)+(in_buffer[94]<<6)+(in_buffer[94]<<9))-(0+(in_buffer[95]<<2)+(in_buffer[95]<<4)+(in_buffer[95]<<8)+(in_buffer[95]<<11))-(0+(in_buffer[96]<<4)-(in_buffer[96]<<7)+(in_buffer[96]<<12))+(0-(in_buffer[97]<<1)-(in_buffer[97]<<3)+(in_buffer[97]<<6)+(in_buffer[97]<<12))+(0+(in_buffer[98]<<4)+(in_buffer[98]<<5)+(in_buffer[98]<<8)+(in_buffer[98]<<10))-(0-(in_buffer[99]<<4)+(in_buffer[99]<<9)+(in_buffer[99]<<11)+(in_buffer[99]<<12))+(0+(in_buffer[100]<<0)+(in_buffer[100]<<2)-(in_buffer[100]<<4)-(in_buffer[100]<<7)+(in_buffer[100]<<11))-(0+(in_buffer[101]<<0)+(in_buffer[101]<<1)+(in_buffer[101]<<4)+(in_buffer[101]<<8)+(in_buffer[101]<<10)+(in_buffer[101]<<12))+(0+(in_buffer[102]<<2)+(in_buffer[102]<<3)+(in_buffer[102]<<6)+(in_buffer[102]<<8))+(0+(in_buffer[103]<<0)-(in_buffer[103]<<2)+(in_buffer[103]<<6)-(in_buffer[103]<<8)+(in_buffer[103]<<12))+(0-(in_buffer[104]<<1)-(in_buffer[104]<<3)+(in_buffer[104]<<6)+(in_buffer[104]<<12))+(0-(in_buffer[105]<<2)+(in_buffer[105]<<7)+(in_buffer[105]<<9)+(in_buffer[105]<<10))+(0-(in_buffer[106]<<0)+(in_buffer[106]<<3)-(in_buffer[106]<<5)+(in_buffer[106]<<7)+(in_buffer[106]<<8)+(in_buffer[106]<<11))-(0+(in_buffer[107]<<6)+(in_buffer[107]<<7)+(in_buffer[107]<<10)+(in_buffer[107]<<12))+(0-(in_buffer[108]<<0)+(in_buffer[108]<<3)+(in_buffer[108]<<4)+(in_buffer[108]<<7)-(in_buffer[108]<<9)+(in_buffer[108]<<12))+(0+(in_buffer[109]<<0)-(in_buffer[109]<<2)-(in_buffer[109]<<5)+(in_buffer[109]<<8)+(in_buffer[109]<<10))-(0+(in_buffer[110]<<1)+(in_buffer[110]<<2)-(in_buffer[110]<<8)+(in_buffer[110]<<10)+(in_buffer[110]<<11))+(0-(in_buffer[111]<<0)+(in_buffer[111]<<5)+(in_buffer[111]<<6)-(in_buffer[111]<<9)+(in_buffer[111]<<11)+(in_buffer[111]<<12))+(0-(in_buffer[112]<<1)+(in_buffer[112]<<5)-(in_buffer[112]<<7)-(in_buffer[112]<<9)+(in_buffer[112]<<12))+(0+(in_buffer[113]<<1)+(in_buffer[113]<<2)-(in_buffer[113]<<6)+(in_buffer[113]<<13))-(0+(in_buffer[114]<<1)+(in_buffer[114]<<2)+(in_buffer[114]<<5)+(in_buffer[114]<<7))-(0-(in_buffer[115]<<3)+(in_buffer[115]<<8)+(in_buffer[115]<<10)+(in_buffer[115]<<11))-(0+(in_buffer[116]<<1)+(in_buffer[116]<<7)+(in_buffer[116]<<8)+(in_buffer[116]<<12))+(0-(in_buffer[117]<<2)-(in_buffer[117]<<5)+(in_buffer[117]<<8)+(in_buffer[117]<<12))+(0+(in_buffer[118]<<1)+(in_buffer[118]<<5)-(in_buffer[118]<<8)+(in_buffer[118]<<11))+(0+(in_buffer[119]<<0)+(in_buffer[119]<<3)+(in_buffer[119]<<5)+(in_buffer[119]<<9)+(in_buffer[119]<<10))-(0-(in_buffer[120]<<1)+(in_buffer[120]<<3)+(in_buffer[120]<<4)+(in_buffer[120]<<7)+(in_buffer[120]<<9)+(in_buffer[120]<<11)+(in_buffer[120]<<12));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight21;
assign in_buffer_weight21=0-(0+(in_buffer[0]<<1)+(in_buffer[0]<<2)+(in_buffer[0]<<7)+(in_buffer[0]<<10)+(in_buffer[0]<<12)+(in_buffer[0]<<13))-(0+(in_buffer[1]<<3)-(in_buffer[1]<<6)-(in_buffer[1]<<8)-(in_buffer[1]<<10)+(in_buffer[1]<<13)+(in_buffer[1]<<14))-(0+(in_buffer[2]<<1)+(in_buffer[2]<<4)+(in_buffer[2]<<7)+(in_buffer[2]<<9)+(in_buffer[2]<<11)+(in_buffer[2]<<14))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<2)+(in_buffer[3]<<6)+(in_buffer[3]<<9))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<1)+(in_buffer[4]<<4)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<0)+(in_buffer[5]<<4)-(in_buffer[5]<<6)-(in_buffer[5]<<8)+(in_buffer[5]<<11))+(0+(in_buffer[6]<<1)+(in_buffer[6]<<2)-(in_buffer[6]<<8)+(in_buffer[6]<<10)+(in_buffer[6]<<11))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<2)+(in_buffer[7]<<4)-(in_buffer[7]<<6)+(in_buffer[7]<<9)+(in_buffer[7]<<12))-(0+(in_buffer[8]<<2)-(in_buffer[8]<<6)-(in_buffer[8]<<11)+(in_buffer[8]<<14))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<1)+(in_buffer[9]<<4)+(in_buffer[9]<<8)+(in_buffer[9]<<10)+(in_buffer[9]<<12))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<5)+(in_buffer[10]<<7)+(in_buffer[10]<<10)+(in_buffer[10]<<11))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3)+(in_buffer[11]<<6)+(in_buffer[11]<<8)+(in_buffer[11]<<10)+(in_buffer[11]<<11))-(0-(in_buffer[12]<<0)-(in_buffer[12]<<3)+(in_buffer[12]<<8)+(in_buffer[12]<<11)+(in_buffer[12]<<12))-(0+(in_buffer[13]<<2)+(in_buffer[13]<<4)+(in_buffer[13]<<8)+(in_buffer[13]<<11))+(0-(in_buffer[14]<<0)-(in_buffer[14]<<2)-(in_buffer[14]<<4)+(in_buffer[14]<<8)+(in_buffer[14]<<9))-(0+(in_buffer[15]<<3)+(in_buffer[15]<<4)+(in_buffer[15]<<7)+(in_buffer[15]<<9))-(0+(in_buffer[16]<<4)+(in_buffer[16]<<5)+(in_buffer[16]<<8)+(in_buffer[16]<<10))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4)+(in_buffer[17]<<6))-(0+(in_buffer[19]<<0)+(in_buffer[19]<<1)-(in_buffer[19]<<7)+(in_buffer[19]<<9)+(in_buffer[19]<<10))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<6)+(in_buffer[20]<<9))+(0-(in_buffer[21]<<1)+(in_buffer[21]<<11)+(in_buffer[21]<<12))-(0-(in_buffer[22]<<1)+(in_buffer[22]<<3)+(in_buffer[22]<<4)+(in_buffer[22]<<7)+(in_buffer[22]<<9)+(in_buffer[22]<<11)+(in_buffer[22]<<12))-(0+(in_buffer[23]<<5)+(in_buffer[23]<<6)+(in_buffer[23]<<9)+(in_buffer[23]<<11))+(0+(in_buffer[24]<<1)+(in_buffer[24]<<3)-(in_buffer[24]<<5)-(in_buffer[24]<<8)+(in_buffer[24]<<12))+(0+(in_buffer[26]<<2)-(in_buffer[26]<<5)+(in_buffer[26]<<10))-(0+(in_buffer[27]<<5)+(in_buffer[27]<<6)+(in_buffer[27]<<9)+(in_buffer[27]<<11))+(0+(in_buffer[28]<<4)+(in_buffer[28]<<5)+(in_buffer[28]<<8)+(in_buffer[28]<<10))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<3)+(in_buffer[29]<<6)+(in_buffer[29]<<10))+(0-(in_buffer[30]<<0)+(in_buffer[30]<<3)-(in_buffer[30]<<6)+(in_buffer[30]<<10)+(in_buffer[30]<<12))+(0-(in_buffer[31]<<1)+(in_buffer[31]<<5)-(in_buffer[31]<<7)-(in_buffer[31]<<9)+(in_buffer[31]<<12))+(0+(in_buffer[32]<<0)+(in_buffer[32]<<2)+(in_buffer[32]<<5)+(in_buffer[32]<<7)+(in_buffer[32]<<10)+(in_buffer[32]<<11))-(0+(in_buffer[33]<<1)-(in_buffer[33]<<3)+(in_buffer[33]<<7)-(in_buffer[33]<<9)+(in_buffer[33]<<13))-(0+(in_buffer[34]<<0)+(in_buffer[34]<<1)-(in_buffer[34]<<5)+(in_buffer[34]<<12))+(0+(in_buffer[35]<<0)+(in_buffer[35]<<1)+(in_buffer[35]<<4)+(in_buffer[35]<<6))-(0+(in_buffer[36]<<1)+(in_buffer[36]<<3)+(in_buffer[36]<<5)-(in_buffer[36]<<7)+(in_buffer[36]<<10)+(in_buffer[36]<<13))-(0+(in_buffer[37]<<0)+(in_buffer[37]<<2)+(in_buffer[37]<<6)+(in_buffer[37]<<9))-(0-(in_buffer[38]<<0)+(in_buffer[38]<<3)+(in_buffer[38]<<4)+(in_buffer[38]<<7)-(in_buffer[38]<<9)+(in_buffer[38]<<12))-(0+(in_buffer[39]<<0)+(in_buffer[39]<<2)+(in_buffer[39]<<3)+(in_buffer[39]<<9)+(in_buffer[39]<<11))-(0+(in_buffer[40]<<3)+(in_buffer[40]<<7)-(in_buffer[40]<<10)+(in_buffer[40]<<13))-(0+(in_buffer[41]<<2)+(in_buffer[41]<<4)+(in_buffer[41]<<8)+(in_buffer[41]<<11))+(0+(in_buffer[42]<<0)+(in_buffer[42]<<4)-(in_buffer[42]<<7)+(in_buffer[42]<<10))+(0+(in_buffer[43]<<0)+(in_buffer[43]<<1)-(in_buffer[43]<<4)-(in_buffer[43]<<6)-(in_buffer[43]<<8)+(in_buffer[43]<<10)+(in_buffer[43]<<11))-(0+(in_buffer[44]<<0)+(in_buffer[44]<<1)-(in_buffer[44]<<5)+(in_buffer[44]<<12))-(0-(in_buffer[45]<<0)+(in_buffer[45]<<10)+(in_buffer[45]<<11))+(0-(in_buffer[46]<<2)+(in_buffer[46]<<7)+(in_buffer[46]<<9)+(in_buffer[46]<<10))-(0+(in_buffer[47]<<0)+(in_buffer[47]<<4)+(in_buffer[47]<<6)+(in_buffer[47]<<11)+(in_buffer[47]<<12))-(0+(in_buffer[48]<<1)+(in_buffer[48]<<2)+(in_buffer[48]<<5)+(in_buffer[48]<<7))-(0+(in_buffer[49]<<0)+(in_buffer[49]<<1)-(in_buffer[49]<<4)-(in_buffer[49]<<6)-(in_buffer[49]<<8)+(in_buffer[49]<<10)+(in_buffer[49]<<11))-(0+(in_buffer[50]<<1)-(in_buffer[50]<<4)+(in_buffer[50]<<9))-(0+(in_buffer[51]<<3)+(in_buffer[51]<<5)+(in_buffer[51]<<9)+(in_buffer[51]<<12))-(0+(in_buffer[52]<<1)+(in_buffer[52]<<2)+(in_buffer[52]<<5)+(in_buffer[52]<<7))+(0+(in_buffer[53]<<0)-(in_buffer[53]<<3)+(in_buffer[53]<<8))+(0+(in_buffer[54]<<0)-(in_buffer[54]<<2)-(in_buffer[54]<<4)+(in_buffer[54]<<7)+(in_buffer[54]<<10)+(in_buffer[54]<<12))+(0-(in_buffer[55]<<3)-(in_buffer[55]<<5)-(in_buffer[55]<<7)+(in_buffer[55]<<11)+(in_buffer[55]<<12))+(0+(in_buffer[56]<<0)+(in_buffer[56]<<3)+(in_buffer[56]<<5)+(in_buffer[56]<<9)+(in_buffer[56]<<10))+(0+(in_buffer[57]<<0)+(in_buffer[57]<<3)+(in_buffer[57]<<5)+(in_buffer[57]<<9)+(in_buffer[57]<<10))+(0+(in_buffer[58]<<1)+(in_buffer[58]<<3)+(in_buffer[58]<<7)+(in_buffer[58]<<10))+(0+(in_buffer[59]<<4)+(in_buffer[59]<<5)+(in_buffer[59]<<8)+(in_buffer[59]<<10))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<6)+(in_buffer[60]<<7)+(in_buffer[60]<<11))-(0-(in_buffer[61]<<0)+(in_buffer[61]<<5)+(in_buffer[61]<<7)+(in_buffer[61]<<8))+(0-(in_buffer[62]<<0)+(in_buffer[62]<<3)-(in_buffer[62]<<5)+(in_buffer[62]<<7)+(in_buffer[62]<<8)+(in_buffer[62]<<11))+(0-(in_buffer[63]<<1)+(in_buffer[63]<<4)-(in_buffer[63]<<6)+(in_buffer[63]<<8)+(in_buffer[63]<<9)+(in_buffer[63]<<12))+(0-(in_buffer[65]<<1)-(in_buffer[65]<<4)+(in_buffer[65]<<7)+(in_buffer[65]<<11))+(0+(in_buffer[66]<<0)-(in_buffer[66]<<4)-(in_buffer[66]<<6)+(in_buffer[66]<<8)+(in_buffer[66]<<9)+(in_buffer[66]<<13))-(0+(in_buffer[67]<<0)+(in_buffer[67]<<3)+(in_buffer[67]<<5)+(in_buffer[67]<<9)+(in_buffer[67]<<10))-(0-(in_buffer[68]<<0)+(in_buffer[68]<<5)+(in_buffer[68]<<7)+(in_buffer[68]<<8))+(0-(in_buffer[69]<<0)+(in_buffer[69]<<2)+(in_buffer[69]<<3)+(in_buffer[69]<<6)+(in_buffer[69]<<8)+(in_buffer[69]<<10)+(in_buffer[69]<<11))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<3)+(in_buffer[70]<<5)+(in_buffer[70]<<9)+(in_buffer[70]<<10))+(0+(in_buffer[71]<<0)+(in_buffer[71]<<2)-(in_buffer[71]<<4)-(in_buffer[71]<<7)+(in_buffer[71]<<11))+(0+(in_buffer[72]<<1)+(in_buffer[72]<<3)+(in_buffer[72]<<7)+(in_buffer[72]<<10))+(0-(in_buffer[73]<<0)+(in_buffer[73]<<2)+(in_buffer[73]<<3)+(in_buffer[73]<<6)+(in_buffer[73]<<8)+(in_buffer[73]<<10)+(in_buffer[73]<<11))+(0-(in_buffer[74]<<0)+(in_buffer[74]<<3)-(in_buffer[74]<<5)+(in_buffer[74]<<7)+(in_buffer[74]<<8)+(in_buffer[74]<<11))-(0-(in_buffer[75]<<0)+(in_buffer[75]<<5)+(in_buffer[75]<<7)+(in_buffer[75]<<8))+(0+(in_buffer[76]<<0)+(in_buffer[76]<<2)+(in_buffer[76]<<4)-(in_buffer[76]<<6)+(in_buffer[76]<<9)+(in_buffer[76]<<12))+(0+(in_buffer[77]<<1)+(in_buffer[77]<<4)+(in_buffer[77]<<6)+(in_buffer[77]<<10)+(in_buffer[77]<<11))-(0+(in_buffer[78]<<1)+(in_buffer[78]<<2)-(in_buffer[78]<<8)+(in_buffer[78]<<10)+(in_buffer[78]<<11))+(0+(in_buffer[79]<<2)-(in_buffer[79]<<5)+(in_buffer[79]<<10))+(0+(in_buffer[80]<<3)+(in_buffer[80]<<5)+(in_buffer[80]<<9)+(in_buffer[80]<<12))+(0+(in_buffer[81]<<0)-(in_buffer[81]<<4)-(in_buffer[81]<<9)+(in_buffer[81]<<12))+(0+(in_buffer[82]<<0)-(in_buffer[82]<<2)-(in_buffer[82]<<4)+(in_buffer[82]<<7)+(in_buffer[82]<<10)+(in_buffer[82]<<12))+(0+(in_buffer[83]<<1)+(in_buffer[83]<<3)+(in_buffer[83]<<7)+(in_buffer[83]<<10))+(0+(in_buffer[84]<<0)-(in_buffer[84]<<3)-(in_buffer[84]<<5)-(in_buffer[84]<<7)+(in_buffer[84]<<10)+(in_buffer[84]<<11))+(0-(in_buffer[85]<<1)-(in_buffer[85]<<4)+(in_buffer[85]<<7)+(in_buffer[85]<<11))-(0-(in_buffer[86]<<1)-(in_buffer[86]<<3)-(in_buffer[86]<<5)+(in_buffer[86]<<9)+(in_buffer[86]<<10))-(0-(in_buffer[87]<<1)-(in_buffer[87]<<3)-(in_buffer[87]<<5)+(in_buffer[87]<<9)+(in_buffer[87]<<10))-(0+(in_buffer[88]<<0)+(in_buffer[88]<<1)+(in_buffer[88]<<4)+(in_buffer[88]<<6))+(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)+(in_buffer[89]<<5)+(in_buffer[89]<<11))+(0+(in_buffer[90]<<0)-(in_buffer[90]<<3)+(in_buffer[90]<<8))-(0+(in_buffer[91]<<3)+(in_buffer[91]<<4)+(in_buffer[91]<<7)+(in_buffer[91]<<9))+(0+(in_buffer[92]<<5)+(in_buffer[92]<<6)+(in_buffer[92]<<9)+(in_buffer[92]<<11))+(0+(in_buffer[93]<<3)-(in_buffer[93]<<6)+(in_buffer[93]<<11))+(0+(in_buffer[94]<<4)+(in_buffer[94]<<5)+(in_buffer[94]<<8)+(in_buffer[94]<<10))-(0-(in_buffer[95]<<1)-(in_buffer[95]<<4)+(in_buffer[95]<<7)+(in_buffer[95]<<11))-(0+(in_buffer[96]<<0)+(in_buffer[96]<<6)+(in_buffer[96]<<7)+(in_buffer[96]<<11))+(0-(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<5)+(in_buffer[97]<<11))-(0+(in_buffer[98]<<1)+(in_buffer[98]<<2)-(in_buffer[98]<<8)+(in_buffer[98]<<10)+(in_buffer[98]<<11))-(0-(in_buffer[99]<<0)-(in_buffer[99]<<2)+(in_buffer[99]<<7)+(in_buffer[99]<<9)+(in_buffer[99]<<12))+(0-(in_buffer[100]<<4)+(in_buffer[100]<<9)+(in_buffer[100]<<11)+(in_buffer[100]<<12))-(0+(in_buffer[101]<<2)+(in_buffer[101]<<4)+(in_buffer[101]<<8)+(in_buffer[101]<<11))-(0+(in_buffer[102]<<2)+(in_buffer[102]<<3)+(in_buffer[102]<<6)+(in_buffer[102]<<8))+(0+(in_buffer[103]<<1)+(in_buffer[103]<<7)+(in_buffer[103]<<8)+(in_buffer[103]<<12))+(0+(in_buffer[104]<<0)+(in_buffer[104]<<4)-(in_buffer[104]<<7)+(in_buffer[104]<<10))+(0+(in_buffer[105]<<0)+(in_buffer[105]<<2)+(in_buffer[105]<<3)+(in_buffer[105]<<9)+(in_buffer[105]<<11))-(0+(in_buffer[106]<<1)+(in_buffer[106]<<2)+(in_buffer[106]<<5)+(in_buffer[106]<<7))-(0-(in_buffer[107]<<1)-(in_buffer[107]<<3)-(in_buffer[107]<<5)+(in_buffer[107]<<9)+(in_buffer[107]<<10))+(0+(in_buffer[108]<<1)+(in_buffer[108]<<7)+(in_buffer[108]<<8)+(in_buffer[108]<<12))-(0+(in_buffer[109]<<1)+(in_buffer[109]<<5)-(in_buffer[109]<<8)+(in_buffer[109]<<11))-(0+(in_buffer[110]<<0)+(in_buffer[110]<<2)+(in_buffer[110]<<4)-(in_buffer[110]<<6)+(in_buffer[110]<<9)+(in_buffer[110]<<12))+(0+(in_buffer[111]<<2)+(in_buffer[111]<<6)-(in_buffer[111]<<9)+(in_buffer[111]<<12))+(0+(in_buffer[112]<<2)+(in_buffer[112]<<3)+(in_buffer[112]<<6)+(in_buffer[112]<<8))+(0+(in_buffer[113]<<4)+(in_buffer[113]<<6)+(in_buffer[113]<<10)+(in_buffer[113]<<13))-(0-(in_buffer[114]<<0)-(in_buffer[114]<<2)+(in_buffer[114]<<5)+(in_buffer[114]<<11))-(0+(in_buffer[115]<<4)-(in_buffer[115]<<7)+(in_buffer[115]<<12))-(0+(in_buffer[116]<<3)+(in_buffer[116]<<5)+(in_buffer[116]<<9)+(in_buffer[116]<<12))+(0+(in_buffer[117]<<0)-(in_buffer[117]<<2)+(in_buffer[117]<<5)+(in_buffer[117]<<7)+(in_buffer[117]<<8)+(in_buffer[117]<<11)+(in_buffer[117]<<12))+(0-(in_buffer[118]<<0)+(in_buffer[118]<<5)+(in_buffer[118]<<7)+(in_buffer[118]<<8))+(0+(in_buffer[119]<<0)+(in_buffer[119]<<2)+(in_buffer[119]<<5)+(in_buffer[119]<<7)+(in_buffer[119]<<10)+(in_buffer[119]<<11))+(0+(in_buffer[120]<<3)+(in_buffer[120]<<4)+(in_buffer[120]<<7)+(in_buffer[120]<<9));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight22;
assign in_buffer_weight22=0+(0+(in_buffer[1]<<2)+(in_buffer[1]<<3)+(in_buffer[1]<<6)+(in_buffer[1]<<8))+(0-(in_buffer[3]<<0)+(in_buffer[3]<<5)+(in_buffer[3]<<7)+(in_buffer[3]<<8))+(0-(in_buffer[4]<<0)-(in_buffer[4]<<2)-(in_buffer[4]<<4)+(in_buffer[4]<<8)+(in_buffer[4]<<9))-(0+(in_buffer[5]<<0)-(in_buffer[5]<<3)+(in_buffer[5]<<8))-(0+(in_buffer[6]<<1)+(in_buffer[6]<<2)+(in_buffer[6]<<5)+(in_buffer[6]<<7))-(0+(in_buffer[7]<<1)-(in_buffer[7]<<4)+(in_buffer[7]<<9))+(0+(in_buffer[9]<<2)+(in_buffer[9]<<3)+(in_buffer[9]<<6)+(in_buffer[9]<<8))-(0+(in_buffer[11]<<3)+(in_buffer[11]<<4)+(in_buffer[11]<<7)+(in_buffer[11]<<9))+(0-(in_buffer[12]<<1)+(in_buffer[12]<<6)+(in_buffer[12]<<8)+(in_buffer[12]<<9))-(0+(in_buffer[13]<<2)+(in_buffer[13]<<3)+(in_buffer[13]<<6)+(in_buffer[13]<<8))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<1)+(in_buffer[15]<<4)+(in_buffer[15]<<6))-(0+(in_buffer[16]<<1)-(in_buffer[16]<<4)+(in_buffer[16]<<9))-(0+(in_buffer[17]<<0)-(in_buffer[17]<<3)+(in_buffer[17]<<8))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<6))-(0+(in_buffer[19]<<1)-(in_buffer[19]<<4)+(in_buffer[19]<<9))-(0-(in_buffer[20]<<0)-(in_buffer[20]<<3)+(in_buffer[20]<<6)+(in_buffer[20]<<10))-(0+(in_buffer[21]<<1)+(in_buffer[21]<<2)+(in_buffer[21]<<5)+(in_buffer[21]<<7))+(0-(in_buffer[23]<<0)-(in_buffer[23]<<2)-(in_buffer[23]<<4)+(in_buffer[23]<<8)+(in_buffer[23]<<9))+(0+(in_buffer[24]<<1)-(in_buffer[24]<<4)+(in_buffer[24]<<9))-(0+(in_buffer[25]<<2)+(in_buffer[25]<<3)+(in_buffer[25]<<6)+(in_buffer[25]<<8))-(0-(in_buffer[26]<<0)-(in_buffer[26]<<2)-(in_buffer[26]<<4)+(in_buffer[26]<<8)+(in_buffer[26]<<9))-(0+(in_buffer[27]<<1)+(in_buffer[27]<<2)+(in_buffer[27]<<5)+(in_buffer[27]<<7))+(0+(in_buffer[28]<<0)-(in_buffer[28]<<3)+(in_buffer[28]<<8))-(0-(in_buffer[29]<<0)-(in_buffer[29]<<3)+(in_buffer[29]<<6)+(in_buffer[29]<<10))-(0+(in_buffer[30]<<0)+(in_buffer[30]<<4)-(in_buffer[30]<<7)+(in_buffer[30]<<10))+(0+(in_buffer[31]<<0)+(in_buffer[31]<<1)+(in_buffer[31]<<4)+(in_buffer[31]<<6))+(0+(in_buffer[32]<<1)-(in_buffer[32]<<4)+(in_buffer[32]<<9))+(0+(in_buffer[35]<<0)+(in_buffer[35]<<4)-(in_buffer[35]<<7)+(in_buffer[35]<<10))-(0+(in_buffer[36]<<0)+(in_buffer[36]<<1)+(in_buffer[36]<<4)+(in_buffer[36]<<6))-(0-(in_buffer[37]<<0)+(in_buffer[37]<<5)+(in_buffer[37]<<7)+(in_buffer[37]<<8))+(0+(in_buffer[38]<<0)-(in_buffer[38]<<3)+(in_buffer[38]<<8))-(0+(in_buffer[39]<<0)+(in_buffer[39]<<2)+(in_buffer[39]<<6)+(in_buffer[39]<<9))-(0+(in_buffer[40]<<0)+(in_buffer[40]<<4)-(in_buffer[40]<<7)+(in_buffer[40]<<10))-(0-(in_buffer[41]<<1)+(in_buffer[41]<<6)+(in_buffer[41]<<8)+(in_buffer[41]<<9))+(0+(in_buffer[44]<<1)-(in_buffer[44]<<4)+(in_buffer[44]<<9))+(0+(in_buffer[45]<<1)+(in_buffer[45]<<2)+(in_buffer[45]<<5)+(in_buffer[45]<<7))+(0+(in_buffer[46]<<0)-(in_buffer[46]<<3)+(in_buffer[46]<<8))+(0+(in_buffer[47]<<2)+(in_buffer[47]<<3)+(in_buffer[47]<<6)+(in_buffer[47]<<8))-(0+(in_buffer[48]<<0)+(in_buffer[48]<<2)+(in_buffer[48]<<6)+(in_buffer[48]<<9))-(0+(in_buffer[49]<<0)-(in_buffer[49]<<3)+(in_buffer[49]<<8))-(0-(in_buffer[50]<<1)+(in_buffer[50]<<6)+(in_buffer[50]<<8)+(in_buffer[50]<<9))-(0+(in_buffer[51]<<0)+(in_buffer[51]<<2)+(in_buffer[51]<<6)+(in_buffer[51]<<9))-(0+(in_buffer[52]<<0)+(in_buffer[52]<<2)+(in_buffer[52]<<6)+(in_buffer[52]<<9))-(0+(in_buffer[54]<<1)-(in_buffer[54]<<4)+(in_buffer[54]<<9))+(0+(in_buffer[55]<<0)-(in_buffer[55]<<3)+(in_buffer[55]<<8))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<6)+(in_buffer[56]<<9))-(0-(in_buffer[57]<<0)-(in_buffer[57]<<2)-(in_buffer[57]<<4)+(in_buffer[57]<<8)+(in_buffer[57]<<9))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)+(in_buffer[58]<<6)+(in_buffer[58]<<9))-(0+(in_buffer[59]<<2)-(in_buffer[59]<<5)+(in_buffer[59]<<10))-(0-(in_buffer[60]<<0)-(in_buffer[60]<<2)-(in_buffer[60]<<4)+(in_buffer[60]<<8)+(in_buffer[60]<<9))-(0+(in_buffer[61]<<0)+(in_buffer[61]<<1)+(in_buffer[61]<<4)+(in_buffer[61]<<6))-(0+(in_buffer[62]<<0)+(in_buffer[62]<<4)-(in_buffer[62]<<7)+(in_buffer[62]<<10))+(0+(in_buffer[64]<<2)+(in_buffer[64]<<3)+(in_buffer[64]<<6)+(in_buffer[64]<<8))-(0+(in_buffer[65]<<0)+(in_buffer[65]<<2)+(in_buffer[65]<<6)+(in_buffer[65]<<9))+(0+(in_buffer[66]<<3)+(in_buffer[66]<<4)+(in_buffer[66]<<7)+(in_buffer[66]<<9))+(0+(in_buffer[67]<<0)+(in_buffer[67]<<1)+(in_buffer[67]<<4)+(in_buffer[67]<<6))-(0+(in_buffer[68]<<3)+(in_buffer[68]<<4)+(in_buffer[68]<<7)+(in_buffer[68]<<9))-(0+(in_buffer[69]<<0)+(in_buffer[69]<<4)-(in_buffer[69]<<7)+(in_buffer[69]<<10))+(0+(in_buffer[70]<<1)-(in_buffer[70]<<4)+(in_buffer[70]<<9))-(0+(in_buffer[71]<<2)+(in_buffer[71]<<3)+(in_buffer[71]<<6)+(in_buffer[71]<<8))+(0+(in_buffer[72]<<2)+(in_buffer[72]<<3)+(in_buffer[72]<<6)+(in_buffer[72]<<8))-(0+(in_buffer[73]<<0)-(in_buffer[73]<<3)+(in_buffer[73]<<8))-(0+(in_buffer[74]<<0)-(in_buffer[74]<<3)+(in_buffer[74]<<8))-(0+(in_buffer[75]<<2)+(in_buffer[75]<<3)+(in_buffer[75]<<6)+(in_buffer[75]<<8))-(0+(in_buffer[76]<<1)-(in_buffer[76]<<4)+(in_buffer[76]<<9))-(0+(in_buffer[77]<<0)-(in_buffer[77]<<3)+(in_buffer[77]<<8))-(0-(in_buffer[78]<<0)+(in_buffer[78]<<5)+(in_buffer[78]<<7)+(in_buffer[78]<<8))+(0+(in_buffer[79]<<0)-(in_buffer[79]<<3)+(in_buffer[79]<<8))+(0+(in_buffer[80]<<0)-(in_buffer[80]<<3)+(in_buffer[80]<<8))-(0+(in_buffer[81]<<0)-(in_buffer[81]<<3)+(in_buffer[81]<<8))+(0+(in_buffer[82]<<2)+(in_buffer[82]<<3)+(in_buffer[82]<<6)+(in_buffer[82]<<8))+(0+(in_buffer[83]<<1)-(in_buffer[83]<<4)+(in_buffer[83]<<9))-(0-(in_buffer[84]<<1)+(in_buffer[84]<<6)+(in_buffer[84]<<8)+(in_buffer[84]<<9))-(0+(in_buffer[85]<<3)+(in_buffer[85]<<4)+(in_buffer[85]<<7)+(in_buffer[85]<<9))-(0+(in_buffer[86]<<0)+(in_buffer[86]<<1)+(in_buffer[86]<<4)+(in_buffer[86]<<6))+(0+(in_buffer[87]<<2)+(in_buffer[87]<<3)+(in_buffer[87]<<6)+(in_buffer[87]<<8))-(0-(in_buffer[88]<<0)-(in_buffer[88]<<3)+(in_buffer[88]<<6)+(in_buffer[88]<<10))-(0+(in_buffer[90]<<1)+(in_buffer[90]<<3)+(in_buffer[90]<<7)+(in_buffer[90]<<10))-(0+(in_buffer[91]<<0)-(in_buffer[91]<<3)+(in_buffer[91]<<8))-(0+(in_buffer[92]<<3)+(in_buffer[92]<<4)+(in_buffer[92]<<7)+(in_buffer[92]<<9))-(0-(in_buffer[93]<<0)-(in_buffer[93]<<3)+(in_buffer[93]<<6)+(in_buffer[93]<<10))-(0+(in_buffer[94]<<0)+(in_buffer[94]<<2)+(in_buffer[94]<<6)+(in_buffer[94]<<9))-(0+(in_buffer[95]<<2)+(in_buffer[95]<<3)+(in_buffer[95]<<6)+(in_buffer[95]<<8))+(0+(in_buffer[96]<<0)-(in_buffer[96]<<3)+(in_buffer[96]<<8))-(0-(in_buffer[97]<<0)+(in_buffer[97]<<5)+(in_buffer[97]<<7)+(in_buffer[97]<<8))-(0-(in_buffer[98]<<0)-(in_buffer[98]<<3)+(in_buffer[98]<<6)+(in_buffer[98]<<10))-(0-(in_buffer[99]<<0)-(in_buffer[99]<<2)-(in_buffer[99]<<4)+(in_buffer[99]<<8)+(in_buffer[99]<<9))-(0-(in_buffer[100]<<0)-(in_buffer[100]<<3)+(in_buffer[100]<<6)+(in_buffer[100]<<10))+(0+(in_buffer[101]<<1)+(in_buffer[101]<<2)+(in_buffer[101]<<5)+(in_buffer[101]<<7))-(0+(in_buffer[102]<<2)+(in_buffer[102]<<3)+(in_buffer[102]<<6)+(in_buffer[102]<<8))-(0+(in_buffer[103]<<0)+(in_buffer[103]<<1)+(in_buffer[103]<<4)+(in_buffer[103]<<6))-(0-(in_buffer[105]<<0)+(in_buffer[105]<<5)+(in_buffer[105]<<7)+(in_buffer[105]<<8))-(0-(in_buffer[106]<<0)-(in_buffer[106]<<2)-(in_buffer[106]<<4)+(in_buffer[106]<<8)+(in_buffer[106]<<9))-(0-(in_buffer[107]<<1)+(in_buffer[107]<<6)+(in_buffer[107]<<8)+(in_buffer[107]<<9))+(0+(in_buffer[108]<<3)+(in_buffer[108]<<4)+(in_buffer[108]<<7)+(in_buffer[108]<<9))+(0+(in_buffer[109]<<1)-(in_buffer[109]<<4)+(in_buffer[109]<<9))-(0+(in_buffer[110]<<0)+(in_buffer[110]<<2)+(in_buffer[110]<<6)+(in_buffer[110]<<9))+(0+(in_buffer[111]<<0)-(in_buffer[111]<<3)+(in_buffer[111]<<8))+(0+(in_buffer[112]<<0)-(in_buffer[112]<<3)+(in_buffer[112]<<8))+(0-(in_buffer[113]<<0)+(in_buffer[113]<<5)+(in_buffer[113]<<7)+(in_buffer[113]<<8))-(0+(in_buffer[114]<<1)-(in_buffer[114]<<4)+(in_buffer[114]<<9))-(0-(in_buffer[115]<<1)+(in_buffer[115]<<6)+(in_buffer[115]<<8)+(in_buffer[115]<<9))+(0-(in_buffer[116]<<0)+(in_buffer[116]<<5)+(in_buffer[116]<<7)+(in_buffer[116]<<8))+(0+(in_buffer[117]<<0)-(in_buffer[117]<<3)+(in_buffer[117]<<8))-(0-(in_buffer[118]<<0)-(in_buffer[118]<<2)-(in_buffer[118]<<4)+(in_buffer[118]<<8)+(in_buffer[118]<<9))-(0+(in_buffer[119]<<3)+(in_buffer[119]<<4)+(in_buffer[119]<<7)+(in_buffer[119]<<9))-(0+(in_buffer[120]<<0)+(in_buffer[120]<<4)-(in_buffer[120]<<7)+(in_buffer[120]<<10));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight23;
assign in_buffer_weight23=0+(0+(in_buffer[0]<<2)+(in_buffer[0]<<3)+(in_buffer[0]<<6)+(in_buffer[0]<<8))+(0+(in_buffer[1]<<1)-(in_buffer[1]<<4)+(in_buffer[1]<<9))+(0-(in_buffer[2]<<0)-(in_buffer[2]<<2)-(in_buffer[2]<<4)+(in_buffer[2]<<8)+(in_buffer[2]<<9))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<2)+(in_buffer[3]<<6)+(in_buffer[3]<<9))-(0+(in_buffer[4]<<1)-(in_buffer[4]<<4)+(in_buffer[4]<<9))+(0+(in_buffer[5]<<2)+(in_buffer[5]<<3)+(in_buffer[5]<<6)+(in_buffer[5]<<8))-(0-(in_buffer[6]<<0)+(in_buffer[6]<<5)+(in_buffer[6]<<7)+(in_buffer[6]<<8))-(0+(in_buffer[7]<<0)+(in_buffer[7]<<1)+(in_buffer[7]<<4)+(in_buffer[7]<<6))-(0+(in_buffer[8]<<2)+(in_buffer[8]<<3)+(in_buffer[8]<<6)+(in_buffer[8]<<8))-(0+(in_buffer[9]<<1)-(in_buffer[9]<<4)+(in_buffer[9]<<9))+(0+(in_buffer[10]<<3)+(in_buffer[10]<<4)+(in_buffer[10]<<7)+(in_buffer[10]<<9))+(0-(in_buffer[11]<<1)+(in_buffer[11]<<6)+(in_buffer[11]<<8)+(in_buffer[11]<<9))-(0-(in_buffer[12]<<1)+(in_buffer[12]<<6)+(in_buffer[12]<<8)+(in_buffer[12]<<9))+(0+(in_buffer[13]<<0)-(in_buffer[13]<<3)+(in_buffer[13]<<8))-(0-(in_buffer[14]<<0)-(in_buffer[14]<<2)-(in_buffer[14]<<4)+(in_buffer[14]<<8)+(in_buffer[14]<<9))-(0-(in_buffer[15]<<1)+(in_buffer[15]<<6)+(in_buffer[15]<<8)+(in_buffer[15]<<9))-(0+(in_buffer[17]<<1)-(in_buffer[17]<<4)+(in_buffer[17]<<9))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<6)+(in_buffer[18]<<9))-(0+(in_buffer[19]<<1)-(in_buffer[19]<<4)+(in_buffer[19]<<9))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<2)+(in_buffer[20]<<5)+(in_buffer[20]<<7))+(0+(in_buffer[21]<<0)-(in_buffer[21]<<3)+(in_buffer[21]<<8))+(0+(in_buffer[22]<<2)+(in_buffer[22]<<3)+(in_buffer[22]<<6)+(in_buffer[22]<<8))+(0+(in_buffer[23]<<1)-(in_buffer[23]<<4)+(in_buffer[23]<<9))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<1)+(in_buffer[24]<<4)+(in_buffer[24]<<6))-(0+(in_buffer[25]<<2)+(in_buffer[25]<<3)+(in_buffer[25]<<6)+(in_buffer[25]<<8))+(0+(in_buffer[26]<<0)-(in_buffer[26]<<3)+(in_buffer[26]<<8))+(0+(in_buffer[27]<<0)-(in_buffer[27]<<3)+(in_buffer[27]<<8))-(0+(in_buffer[28]<<3)+(in_buffer[28]<<4)+(in_buffer[28]<<7)+(in_buffer[28]<<9))+(0+(in_buffer[29]<<2)+(in_buffer[29]<<3)+(in_buffer[29]<<6)+(in_buffer[29]<<8))-(0+(in_buffer[30]<<1)+(in_buffer[30]<<2)+(in_buffer[30]<<5)+(in_buffer[30]<<7))-(0+(in_buffer[32]<<1)+(in_buffer[32]<<2)+(in_buffer[32]<<5)+(in_buffer[32]<<7))+(0+(in_buffer[33]<<2)+(in_buffer[33]<<3)+(in_buffer[33]<<6)+(in_buffer[33]<<8))+(0-(in_buffer[34]<<0)+(in_buffer[34]<<5)+(in_buffer[34]<<7)+(in_buffer[34]<<8))+(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)-(in_buffer[36]<<4)+(in_buffer[36]<<8)+(in_buffer[36]<<9))+(0+(in_buffer[37]<<0)-(in_buffer[37]<<3)+(in_buffer[37]<<8))+(0+(in_buffer[38]<<0)+(in_buffer[38]<<2)+(in_buffer[38]<<6)+(in_buffer[38]<<9))-(0+(in_buffer[39]<<2)-(in_buffer[39]<<5)+(in_buffer[39]<<10))-(0-(in_buffer[40]<<0)-(in_buffer[40]<<2)-(in_buffer[40]<<4)+(in_buffer[40]<<8)+(in_buffer[40]<<9))+(0-(in_buffer[41]<<1)+(in_buffer[41]<<6)+(in_buffer[41]<<8)+(in_buffer[41]<<9))+(0+(in_buffer[42]<<3)+(in_buffer[42]<<4)+(in_buffer[42]<<7)+(in_buffer[42]<<9))+(0-(in_buffer[43]<<0)+(in_buffer[43]<<5)+(in_buffer[43]<<7)+(in_buffer[43]<<8))+(0+(in_buffer[44]<<0)+(in_buffer[44]<<2)+(in_buffer[44]<<6)+(in_buffer[44]<<9))+(0+(in_buffer[45]<<3)+(in_buffer[45]<<4)+(in_buffer[45]<<7)+(in_buffer[45]<<9))-(0+(in_buffer[46]<<0)+(in_buffer[46]<<4)-(in_buffer[46]<<7)+(in_buffer[46]<<10))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<1)+(in_buffer[47]<<4)+(in_buffer[47]<<6))-(0-(in_buffer[48]<<0)+(in_buffer[48]<<5)+(in_buffer[48]<<7)+(in_buffer[48]<<8))-(0+(in_buffer[49]<<2)+(in_buffer[49]<<3)+(in_buffer[49]<<6)+(in_buffer[49]<<8))-(0+(in_buffer[50]<<0)+(in_buffer[50]<<2)+(in_buffer[50]<<6)+(in_buffer[50]<<9))-(0+(in_buffer[51]<<0)+(in_buffer[51]<<4)-(in_buffer[51]<<7)+(in_buffer[51]<<10))-(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)-(in_buffer[52]<<4)+(in_buffer[52]<<8)+(in_buffer[52]<<9))-(0+(in_buffer[53]<<1)-(in_buffer[53]<<4)+(in_buffer[53]<<9))-(0+(in_buffer[54]<<0)+(in_buffer[54]<<1)+(in_buffer[54]<<4)+(in_buffer[54]<<6))-(0+(in_buffer[55]<<2)+(in_buffer[55]<<3)+(in_buffer[55]<<6)+(in_buffer[55]<<8))+(0+(in_buffer[56]<<1)-(in_buffer[56]<<4)+(in_buffer[56]<<9))+(0-(in_buffer[57]<<0)-(in_buffer[57]<<2)-(in_buffer[57]<<4)+(in_buffer[57]<<8)+(in_buffer[57]<<9))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)+(in_buffer[58]<<6)+(in_buffer[58]<<9))-(0-(in_buffer[59]<<0)-(in_buffer[59]<<2)-(in_buffer[59]<<4)+(in_buffer[59]<<8)+(in_buffer[59]<<9))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<4)-(in_buffer[60]<<7)+(in_buffer[60]<<10))+(0-(in_buffer[61]<<1)+(in_buffer[61]<<6)+(in_buffer[61]<<8)+(in_buffer[61]<<9))+(0+(in_buffer[62]<<0)-(in_buffer[62]<<3)+(in_buffer[62]<<8))+(0-(in_buffer[63]<<0)-(in_buffer[63]<<2)-(in_buffer[63]<<4)+(in_buffer[63]<<8)+(in_buffer[63]<<9))+(0+(in_buffer[64]<<2)+(in_buffer[64]<<3)+(in_buffer[64]<<6)+(in_buffer[64]<<8))+(0+(in_buffer[65]<<1)-(in_buffer[65]<<4)+(in_buffer[65]<<9))-(0+(in_buffer[66]<<0)+(in_buffer[66]<<2)+(in_buffer[66]<<6)+(in_buffer[66]<<9))-(0+(in_buffer[67]<<3)+(in_buffer[67]<<4)+(in_buffer[67]<<7)+(in_buffer[67]<<9))-(0-(in_buffer[68]<<0)-(in_buffer[68]<<2)-(in_buffer[68]<<4)+(in_buffer[68]<<8)+(in_buffer[68]<<9))-(0-(in_buffer[69]<<1)+(in_buffer[69]<<6)+(in_buffer[69]<<8)+(in_buffer[69]<<9))+(0+(in_buffer[70]<<2)+(in_buffer[70]<<3)+(in_buffer[70]<<6)+(in_buffer[70]<<8))+(0-(in_buffer[71]<<1)+(in_buffer[71]<<6)+(in_buffer[71]<<8)+(in_buffer[71]<<9))-(0+(in_buffer[72]<<0)+(in_buffer[72]<<4)-(in_buffer[72]<<7)+(in_buffer[72]<<10))+(0+(in_buffer[73]<<3)+(in_buffer[73]<<4)+(in_buffer[73]<<7)+(in_buffer[73]<<9))+(0+(in_buffer[74]<<0)+(in_buffer[74]<<2)+(in_buffer[74]<<6)+(in_buffer[74]<<9))+(0+(in_buffer[75]<<0)-(in_buffer[75]<<3)+(in_buffer[75]<<8))-(0+(in_buffer[76]<<0)+(in_buffer[76]<<4)-(in_buffer[76]<<7)+(in_buffer[76]<<10))-(0+(in_buffer[77]<<1)-(in_buffer[77]<<4)+(in_buffer[77]<<9))+(0+(in_buffer[78]<<0)-(in_buffer[78]<<3)+(in_buffer[78]<<8))-(0-(in_buffer[79]<<0)+(in_buffer[79]<<5)+(in_buffer[79]<<7)+(in_buffer[79]<<8))+(0+(in_buffer[80]<<3)+(in_buffer[80]<<4)+(in_buffer[80]<<7)+(in_buffer[80]<<9))+(0+(in_buffer[81]<<0)+(in_buffer[81]<<1)+(in_buffer[81]<<4)+(in_buffer[81]<<6))-(0+(in_buffer[82]<<1)+(in_buffer[82]<<2)+(in_buffer[82]<<5)+(in_buffer[82]<<7))-(0-(in_buffer[83]<<0)-(in_buffer[83]<<2)-(in_buffer[83]<<4)+(in_buffer[83]<<8)+(in_buffer[83]<<9))+(0+(in_buffer[85]<<0)+(in_buffer[85]<<1)+(in_buffer[85]<<4)+(in_buffer[85]<<6))-(0-(in_buffer[86]<<0)+(in_buffer[86]<<5)+(in_buffer[86]<<7)+(in_buffer[86]<<8))-(0+(in_buffer[87]<<0)-(in_buffer[87]<<3)+(in_buffer[87]<<8))-(0-(in_buffer[88]<<1)+(in_buffer[88]<<6)+(in_buffer[88]<<8)+(in_buffer[88]<<9))+(0+(in_buffer[89]<<2)+(in_buffer[89]<<3)+(in_buffer[89]<<6)+(in_buffer[89]<<8))+(0+(in_buffer[90]<<1)-(in_buffer[90]<<4)+(in_buffer[90]<<9))+(0+(in_buffer[91]<<0)+(in_buffer[91]<<2)+(in_buffer[91]<<6)+(in_buffer[91]<<9))-(0+(in_buffer[92]<<2)+(in_buffer[92]<<3)+(in_buffer[92]<<6)+(in_buffer[92]<<8))-(0+(in_buffer[93]<<0)+(in_buffer[93]<<2)+(in_buffer[93]<<6)+(in_buffer[93]<<9))-(0+(in_buffer[95]<<0)+(in_buffer[95]<<4)-(in_buffer[95]<<7)+(in_buffer[95]<<10))-(0+(in_buffer[96]<<2)-(in_buffer[96]<<5)+(in_buffer[96]<<10))-(0-(in_buffer[97]<<0)+(in_buffer[97]<<5)+(in_buffer[97]<<7)+(in_buffer[97]<<8))-(0+(in_buffer[98]<<0)+(in_buffer[98]<<2)+(in_buffer[98]<<6)+(in_buffer[98]<<9))+(0-(in_buffer[99]<<0)+(in_buffer[99]<<5)+(in_buffer[99]<<7)+(in_buffer[99]<<8))+(0+(in_buffer[100]<<0)-(in_buffer[100]<<3)+(in_buffer[100]<<8))+(0-(in_buffer[101]<<0)+(in_buffer[101]<<5)+(in_buffer[101]<<7)+(in_buffer[101]<<8))+(0+(in_buffer[102]<<1)-(in_buffer[102]<<4)+(in_buffer[102]<<9))-(0+(in_buffer[103]<<0)+(in_buffer[103]<<4)-(in_buffer[103]<<7)+(in_buffer[103]<<10))-(0+(in_buffer[104]<<1)+(in_buffer[104]<<2)+(in_buffer[104]<<5)+(in_buffer[104]<<7))-(0+(in_buffer[105]<<3)+(in_buffer[105]<<4)+(in_buffer[105]<<7)+(in_buffer[105]<<9))-(0-(in_buffer[106]<<0)-(in_buffer[106]<<2)-(in_buffer[106]<<4)+(in_buffer[106]<<8)+(in_buffer[106]<<9))+(0+(in_buffer[107]<<0)-(in_buffer[107]<<3)+(in_buffer[107]<<8))+(0+(in_buffer[108]<<2)+(in_buffer[108]<<3)+(in_buffer[108]<<6)+(in_buffer[108]<<8))+(0+(in_buffer[109]<<0)+(in_buffer[109]<<2)+(in_buffer[109]<<6)+(in_buffer[109]<<9))+(0+(in_buffer[110]<<2)+(in_buffer[110]<<3)+(in_buffer[110]<<6)+(in_buffer[110]<<8))-(0-(in_buffer[111]<<1)+(in_buffer[111]<<6)+(in_buffer[111]<<8)+(in_buffer[111]<<9))-(0-(in_buffer[113]<<1)+(in_buffer[113]<<6)+(in_buffer[113]<<8)+(in_buffer[113]<<9))+(0+(in_buffer[114]<<0)+(in_buffer[114]<<2)+(in_buffer[114]<<6)+(in_buffer[114]<<9))+(0+(in_buffer[115]<<1)+(in_buffer[115]<<2)+(in_buffer[115]<<5)+(in_buffer[115]<<7))+(0+(in_buffer[116]<<3)+(in_buffer[116]<<4)+(in_buffer[116]<<7)+(in_buffer[116]<<9))-(0+(in_buffer[117]<<3)+(in_buffer[117]<<4)+(in_buffer[117]<<7)+(in_buffer[117]<<9))+(0+(in_buffer[118]<<2)+(in_buffer[118]<<3)+(in_buffer[118]<<6)+(in_buffer[118]<<8))+(0-(in_buffer[119]<<0)+(in_buffer[119]<<5)+(in_buffer[119]<<7)+(in_buffer[119]<<8));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight24;
assign in_buffer_weight24=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<10)+(in_buffer[0]<<11))-(0+(in_buffer[1]<<2)+(in_buffer[1]<<5)+(in_buffer[1]<<7)+(in_buffer[1]<<11)+(in_buffer[1]<<12))+(0-(in_buffer[2]<<2)+(in_buffer[2]<<5)-(in_buffer[2]<<7)+(in_buffer[2]<<9)+(in_buffer[2]<<10)+(in_buffer[2]<<13))+(0+(in_buffer[3]<<0)-(in_buffer[3]<<3)-(in_buffer[3]<<6)-(in_buffer[3]<<9)+(in_buffer[3]<<11)+(in_buffer[3]<<12))+(0-(in_buffer[4]<<1)-(in_buffer[4]<<4)+(in_buffer[4]<<7)+(in_buffer[4]<<11))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<3)+(in_buffer[5]<<5)-(in_buffer[5]<<7)+(in_buffer[5]<<10)+(in_buffer[5]<<13))-(0-(in_buffer[6]<<3)+(in_buffer[6]<<8)+(in_buffer[6]<<10)+(in_buffer[6]<<11))+(0+(in_buffer[7]<<0)+(in_buffer[7]<<1)-(in_buffer[7]<<4)-(in_buffer[7]<<6)-(in_buffer[7]<<8)+(in_buffer[7]<<10)+(in_buffer[7]<<11))+(0-(in_buffer[8]<<1)-(in_buffer[8]<<3)+(in_buffer[8]<<8)+(in_buffer[8]<<10)+(in_buffer[8]<<13))-(0+(in_buffer[9]<<1)+(in_buffer[9]<<2)-(in_buffer[9]<<5)-(in_buffer[9]<<7)-(in_buffer[9]<<9)+(in_buffer[9]<<11)+(in_buffer[9]<<12))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<3)-(in_buffer[10]<<7)+(in_buffer[10]<<10)+(in_buffer[10]<<12)+(in_buffer[10]<<13))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<1)-(in_buffer[11]<<4)-(in_buffer[11]<<6)-(in_buffer[11]<<8)+(in_buffer[11]<<10)+(in_buffer[11]<<11))+(0+(in_buffer[12]<<2)+(in_buffer[12]<<4)-(in_buffer[12]<<6)-(in_buffer[12]<<9)+(in_buffer[12]<<13))+(0+(in_buffer[13]<<0)-(in_buffer[13]<<4)-(in_buffer[13]<<9)+(in_buffer[13]<<12))-(0-(in_buffer[14]<<0)+(in_buffer[14]<<10)+(in_buffer[14]<<11))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3)+(in_buffer[15]<<9)+(in_buffer[15]<<11))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<10)+(in_buffer[16]<<11))-(0+(in_buffer[17]<<3)-(in_buffer[17]<<6)+(in_buffer[17]<<11))-(0-(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<7)+(in_buffer[18]<<9)+(in_buffer[18]<<12))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<1)-(in_buffer[19]<<4)-(in_buffer[19]<<6)-(in_buffer[19]<<8)+(in_buffer[19]<<10)+(in_buffer[19]<<11))+(0-(in_buffer[20]<<2)-(in_buffer[20]<<5)+(in_buffer[20]<<8)+(in_buffer[20]<<12))-(0+(in_buffer[21]<<0)-(in_buffer[21]<<2)+(in_buffer[21]<<10)+(in_buffer[21]<<13))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<1)-(in_buffer[22]<<7)+(in_buffer[22]<<9)+(in_buffer[22]<<10))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<2)+(in_buffer[23]<<4)-(in_buffer[23]<<6)+(in_buffer[23]<<9)+(in_buffer[23]<<12))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<2)-(in_buffer[24]<<4)-(in_buffer[24]<<7)+(in_buffer[24]<<11))+(0+(in_buffer[25]<<0)+(in_buffer[25]<<2)-(in_buffer[25]<<4)-(in_buffer[25]<<7)+(in_buffer[25]<<11))-(0-(in_buffer[26]<<0)+(in_buffer[26]<<4)+(in_buffer[26]<<5)+(in_buffer[26]<<8)+(in_buffer[26]<<12))-(0+(in_buffer[27]<<0)+(in_buffer[27]<<1)+(in_buffer[27]<<4)+(in_buffer[27]<<6))-(0+(in_buffer[28]<<0)-(in_buffer[28]<<2)-(in_buffer[28]<<5)+(in_buffer[28]<<8)+(in_buffer[28]<<10))-(0-(in_buffer[29]<<0)+(in_buffer[29]<<5)+(in_buffer[29]<<6)-(in_buffer[29]<<9)+(in_buffer[29]<<11)+(in_buffer[29]<<12))+(0+(in_buffer[30]<<0)-(in_buffer[30]<<3)-(in_buffer[30]<<6)-(in_buffer[30]<<9)+(in_buffer[30]<<11)+(in_buffer[30]<<12))+(0-(in_buffer[31]<<2)-(in_buffer[31]<<5)+(in_buffer[31]<<8)+(in_buffer[31]<<12))-(0-(in_buffer[32]<<1)+(in_buffer[32]<<4)+(in_buffer[32]<<5)+(in_buffer[32]<<8)-(in_buffer[32]<<10)+(in_buffer[32]<<13))-(0+(in_buffer[33]<<0)+(in_buffer[33]<<2)+(in_buffer[33]<<6)+(in_buffer[33]<<9))-(0+(in_buffer[34]<<0)+(in_buffer[34]<<6)+(in_buffer[34]<<7)+(in_buffer[34]<<11))+(0+(in_buffer[35]<<3)-(in_buffer[35]<<6)+(in_buffer[35]<<11))+(0-(in_buffer[36]<<0)-(in_buffer[36]<<2)+(in_buffer[36]<<7)+(in_buffer[36]<<9)+(in_buffer[36]<<12))+(0-(in_buffer[38]<<0)-(in_buffer[38]<<3)+(in_buffer[38]<<8)+(in_buffer[38]<<11)+(in_buffer[38]<<12))-(0+(in_buffer[39]<<5)+(in_buffer[39]<<6)+(in_buffer[39]<<9)+(in_buffer[39]<<11))-(0-(in_buffer[40]<<1)+(in_buffer[40]<<6)+(in_buffer[40]<<8)+(in_buffer[40]<<9))+(0+(in_buffer[41]<<0)+(in_buffer[41]<<2)+(in_buffer[41]<<4)+(in_buffer[41]<<5)-(in_buffer[41]<<10)+(in_buffer[41]<<13))-(0-(in_buffer[42]<<2)-(in_buffer[42]<<5)+(in_buffer[42]<<8)+(in_buffer[42]<<12))+(0+(in_buffer[43]<<1)-(in_buffer[43]<<4)+(in_buffer[43]<<9))-(0-(in_buffer[44]<<1)+(in_buffer[44]<<5)-(in_buffer[44]<<7)-(in_buffer[44]<<9)+(in_buffer[44]<<12))-(0+(in_buffer[45]<<2)+(in_buffer[45]<<6)-(in_buffer[45]<<9)+(in_buffer[45]<<12))+(0-(in_buffer[46]<<1)-(in_buffer[46]<<3)+(in_buffer[46]<<6)+(in_buffer[46]<<12))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<4)-(in_buffer[47]<<7)+(in_buffer[47]<<10))-(0+(in_buffer[48]<<3)+(in_buffer[48]<<5)+(in_buffer[48]<<9)+(in_buffer[48]<<12))+(0+(in_buffer[50]<<0)-(in_buffer[50]<<2)-(in_buffer[50]<<5)+(in_buffer[50]<<8)+(in_buffer[50]<<10))-(0+(in_buffer[51]<<3)+(in_buffer[51]<<4)+(in_buffer[51]<<7)+(in_buffer[51]<<9))+(0-(in_buffer[52]<<1)-(in_buffer[52]<<3)+(in_buffer[52]<<6)+(in_buffer[52]<<12))-(0+(in_buffer[53]<<0)+(in_buffer[53]<<3)+(in_buffer[53]<<5)+(in_buffer[53]<<9)+(in_buffer[53]<<10))-(0-(in_buffer[54]<<1)+(in_buffer[54]<<6)+(in_buffer[54]<<8)+(in_buffer[54]<<9))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<3)+(in_buffer[56]<<7)+(in_buffer[56]<<12))+(0+(in_buffer[57]<<0)+(in_buffer[57]<<1)+(in_buffer[57]<<6)+(in_buffer[57]<<9)+(in_buffer[57]<<11)+(in_buffer[57]<<12))-(0+(in_buffer[58]<<1)+(in_buffer[58]<<5)-(in_buffer[58]<<8)+(in_buffer[58]<<11))+(0-(in_buffer[59]<<0)+(in_buffer[59]<<3)-(in_buffer[59]<<5)+(in_buffer[59]<<7)+(in_buffer[59]<<8)+(in_buffer[59]<<11))+(0-(in_buffer[60]<<1)+(in_buffer[60]<<6)+(in_buffer[60]<<8)+(in_buffer[60]<<9))+(0-(in_buffer[61]<<1)+(in_buffer[61]<<6)+(in_buffer[61]<<8)+(in_buffer[61]<<9))-(0-(in_buffer[62]<<0)+(in_buffer[62]<<4)-(in_buffer[62]<<6)-(in_buffer[62]<<8)+(in_buffer[62]<<11))+(0+(in_buffer[63]<<0)-(in_buffer[63]<<2)-(in_buffer[63]<<5)+(in_buffer[63]<<8)+(in_buffer[63]<<10))-(0+(in_buffer[64]<<0)-(in_buffer[64]<<2)-(in_buffer[64]<<5)+(in_buffer[64]<<8)+(in_buffer[64]<<10))-(0+(in_buffer[65]<<1)+(in_buffer[65]<<3)+(in_buffer[65]<<4)+(in_buffer[65]<<10)+(in_buffer[65]<<12))-(0+(in_buffer[66]<<0)+(in_buffer[66]<<3)+(in_buffer[66]<<7)+(in_buffer[66]<<12))-(0-(in_buffer[67]<<1)-(in_buffer[67]<<3)-(in_buffer[67]<<5)+(in_buffer[67]<<9)+(in_buffer[67]<<10))+(0+(in_buffer[68]<<0)+(in_buffer[68]<<2)+(in_buffer[68]<<3)-(in_buffer[68]<<6)-(in_buffer[68]<<8)+(in_buffer[68]<<13))-(0+(in_buffer[69]<<2)-(in_buffer[69]<<5)+(in_buffer[69]<<10))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<2)+(in_buffer[70]<<6)+(in_buffer[70]<<9))+(0-(in_buffer[71]<<0)+(in_buffer[71]<<4)-(in_buffer[71]<<6)-(in_buffer[71]<<8)+(in_buffer[71]<<11))+(0-(in_buffer[72]<<2)+(in_buffer[72]<<7)+(in_buffer[72]<<9)+(in_buffer[72]<<10))-(0+(in_buffer[73]<<0)+(in_buffer[73]<<2)+(in_buffer[73]<<6)+(in_buffer[73]<<9))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6)-(in_buffer[74]<<8)+(in_buffer[74]<<12))-(0+(in_buffer[75]<<1)+(in_buffer[75]<<2)-(in_buffer[75]<<8)+(in_buffer[75]<<10)+(in_buffer[75]<<11))+(0+(in_buffer[76]<<0)+(in_buffer[76]<<3)+(in_buffer[76]<<5)+(in_buffer[76]<<9)+(in_buffer[76]<<10))+(0+(in_buffer[77]<<1)+(in_buffer[77]<<2)+(in_buffer[77]<<5)+(in_buffer[77]<<7))-(0+(in_buffer[78]<<0)-(in_buffer[78]<<2)-(in_buffer[78]<<5)+(in_buffer[78]<<8)+(in_buffer[78]<<10))+(0-(in_buffer[79]<<1)-(in_buffer[79]<<3)+(in_buffer[79]<<6)+(in_buffer[79]<<12))-(0+(in_buffer[80]<<0)-(in_buffer[80]<<3)-(in_buffer[80]<<5)-(in_buffer[80]<<7)+(in_buffer[80]<<10)+(in_buffer[80]<<11))+(0+(in_buffer[81]<<0)+(in_buffer[81]<<2)-(in_buffer[81]<<4)-(in_buffer[81]<<7)+(in_buffer[81]<<11))+(0-(in_buffer[83]<<0)+(in_buffer[83]<<2)+(in_buffer[83]<<3)+(in_buffer[83]<<6)+(in_buffer[83]<<8)+(in_buffer[83]<<10)+(in_buffer[83]<<11))-(0+(in_buffer[84]<<2)-(in_buffer[84]<<4)-(in_buffer[84]<<7)+(in_buffer[84]<<10)+(in_buffer[84]<<12))+(0+(in_buffer[85]<<1)+(in_buffer[85]<<5)-(in_buffer[85]<<8)+(in_buffer[85]<<11))+(0+(in_buffer[86]<<0)-(in_buffer[86]<<3)-(in_buffer[86]<<5)-(in_buffer[86]<<7)+(in_buffer[86]<<10)+(in_buffer[86]<<11))+(0-(in_buffer[87]<<1)+(in_buffer[87]<<6)+(in_buffer[87]<<8)+(in_buffer[87]<<9))+(0-(in_buffer[88]<<0)+(in_buffer[88]<<10)+(in_buffer[88]<<11))-(0-(in_buffer[89]<<0)-(in_buffer[89]<<2)-(in_buffer[89]<<4)+(in_buffer[89]<<8)+(in_buffer[89]<<9))+(0-(in_buffer[90]<<1)-(in_buffer[90]<<3)+(in_buffer[90]<<6)+(in_buffer[90]<<12))-(0-(in_buffer[91]<<0)+(in_buffer[91]<<5)+(in_buffer[91]<<7)+(in_buffer[91]<<8))+(0-(in_buffer[92]<<0)+(in_buffer[92]<<3)-(in_buffer[92]<<6)+(in_buffer[92]<<10)+(in_buffer[92]<<12))-(0+(in_buffer[93]<<0)+(in_buffer[93]<<4)-(in_buffer[93]<<7)+(in_buffer[93]<<10))-(0+(in_buffer[94]<<4)+(in_buffer[94]<<5)+(in_buffer[94]<<8)+(in_buffer[94]<<10))-(0-(in_buffer[95]<<1)+(in_buffer[95]<<6)+(in_buffer[95]<<7)-(in_buffer[95]<<10)+(in_buffer[95]<<12)+(in_buffer[95]<<13))+(0-(in_buffer[96]<<1)+(in_buffer[96]<<5)-(in_buffer[96]<<7)-(in_buffer[96]<<9)+(in_buffer[96]<<12))+(0-(in_buffer[97]<<2)-(in_buffer[97]<<5)+(in_buffer[97]<<8)+(in_buffer[97]<<12))+(0+(in_buffer[98]<<1)+(in_buffer[98]<<2)+(in_buffer[98]<<5)+(in_buffer[98]<<7))+(0+(in_buffer[99]<<0)+(in_buffer[99]<<2)-(in_buffer[99]<<4)-(in_buffer[99]<<7)+(in_buffer[99]<<11))+(0+(in_buffer[100]<<0)+(in_buffer[100]<<1)+(in_buffer[100]<<4)+(in_buffer[100]<<6))+(0-(in_buffer[101]<<2)+(in_buffer[101]<<7)+(in_buffer[101]<<9)+(in_buffer[101]<<10))-(0-(in_buffer[102]<<1)+(in_buffer[102]<<6)+(in_buffer[102]<<8)+(in_buffer[102]<<9))+(0+(in_buffer[103]<<0)-(in_buffer[103]<<3)-(in_buffer[103]<<5)-(in_buffer[103]<<7)+(in_buffer[103]<<10)+(in_buffer[103]<<11))-(0-(in_buffer[104]<<0)+(in_buffer[104]<<4)-(in_buffer[104]<<6)-(in_buffer[104]<<8)+(in_buffer[104]<<11))+(0-(in_buffer[105]<<0)+(in_buffer[105]<<5)+(in_buffer[105]<<7)+(in_buffer[105]<<8))-(0+(in_buffer[106]<<0)+(in_buffer[106]<<2)-(in_buffer[106]<<8)+(in_buffer[106]<<11)+(in_buffer[106]<<12))+(0-(in_buffer[107]<<0)+(in_buffer[107]<<4)-(in_buffer[107]<<6)-(in_buffer[107]<<8)+(in_buffer[107]<<11))+(0+(in_buffer[108]<<0)-(in_buffer[108]<<2)-(in_buffer[108]<<5)+(in_buffer[108]<<8)+(in_buffer[108]<<10))+(0+(in_buffer[109]<<0)-(in_buffer[109]<<3)-(in_buffer[109]<<5)-(in_buffer[109]<<7)+(in_buffer[109]<<10)+(in_buffer[109]<<11))+(0+(in_buffer[110]<<5)+(in_buffer[110]<<6)+(in_buffer[110]<<9)+(in_buffer[110]<<11))+(0+(in_buffer[111]<<0)+(in_buffer[111]<<1)+(in_buffer[111]<<4)+(in_buffer[111]<<6))+(0-(in_buffer[112]<<0)+(in_buffer[112]<<3)+(in_buffer[112]<<4)+(in_buffer[112]<<7)-(in_buffer[112]<<9)+(in_buffer[112]<<12))-(0+(in_buffer[113]<<0)+(in_buffer[113]<<1)-(in_buffer[113]<<5)+(in_buffer[113]<<12))+(0+(in_buffer[114]<<0)+(in_buffer[114]<<1)+(in_buffer[114]<<4)+(in_buffer[114]<<6))-(0-(in_buffer[115]<<1)+(in_buffer[115]<<3)+(in_buffer[115]<<4)+(in_buffer[115]<<7)+(in_buffer[115]<<9)+(in_buffer[115]<<11)+(in_buffer[115]<<12))+(0+(in_buffer[116]<<1)+(in_buffer[116]<<2)-(in_buffer[116]<<8)+(in_buffer[116]<<10)+(in_buffer[116]<<11))-(0+(in_buffer[117]<<1)-(in_buffer[117]<<3)-(in_buffer[117]<<6)+(in_buffer[117]<<9)+(in_buffer[117]<<11))+(0-(in_buffer[118]<<0)-(in_buffer[118]<<3)+(in_buffer[118]<<8)+(in_buffer[118]<<11)+(in_buffer[118]<<12))+(0+(in_buffer[119]<<0)+(in_buffer[119]<<4)-(in_buffer[119]<<7)+(in_buffer[119]<<10))-(0+(in_buffer[120]<<0)+(in_buffer[120]<<1)+(in_buffer[120]<<4)+(in_buffer[120]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight25;
assign in_buffer_weight25=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<6)+(in_buffer[0]<<7)+(in_buffer[0]<<13))+(0-(in_buffer[1]<<2)-(in_buffer[1]<<4)-(in_buffer[1]<<6)+(in_buffer[1]<<10)+(in_buffer[1]<<11))+(0-(in_buffer[2]<<0)+(in_buffer[2]<<3)-(in_buffer[2]<<5)+(in_buffer[2]<<7)+(in_buffer[2]<<8)+(in_buffer[2]<<11))+(0+(in_buffer[3]<<1)-(in_buffer[3]<<3)-(in_buffer[3]<<6)+(in_buffer[3]<<9)+(in_buffer[3]<<11))-(0-(in_buffer[4]<<0)-(in_buffer[4]<<2)-(in_buffer[4]<<4)+(in_buffer[4]<<7)-(in_buffer[4]<<10)+(in_buffer[4]<<12)+(in_buffer[4]<<13))-(0+(in_buffer[5]<<0)-(in_buffer[5]<<2)-(in_buffer[5]<<4)-(in_buffer[5]<<9)+(in_buffer[5]<<14))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<1)+(in_buffer[6]<<5)+(in_buffer[6]<<7)+(in_buffer[6]<<10)+(in_buffer[6]<<13))-(0+(in_buffer[7]<<2)+(in_buffer[7]<<4)+(in_buffer[7]<<8)+(in_buffer[7]<<11))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<4)-(in_buffer[8]<<6)-(in_buffer[8]<<8)+(in_buffer[8]<<11))+(0+(in_buffer[9]<<2)+(in_buffer[9]<<3)+(in_buffer[9]<<6)+(in_buffer[9]<<8))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)-(in_buffer[10]<<4)-(in_buffer[10]<<6)-(in_buffer[10]<<8)+(in_buffer[10]<<10)+(in_buffer[10]<<11))-(0+(in_buffer[11]<<3)+(in_buffer[11]<<4)+(in_buffer[11]<<7)+(in_buffer[11]<<9))-(0+(in_buffer[12]<<1)-(in_buffer[12]<<3)+(in_buffer[12]<<7)-(in_buffer[12]<<9)+(in_buffer[12]<<13))+(0+(in_buffer[13]<<0)+(in_buffer[13]<<1)+(in_buffer[13]<<4)+(in_buffer[13]<<6))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<5)+(in_buffer[14]<<8)+(in_buffer[14]<<9)+(in_buffer[14]<<12))+(0+(in_buffer[15]<<1)+(in_buffer[15]<<5)-(in_buffer[15]<<8)+(in_buffer[15]<<11))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<5)+(in_buffer[16]<<7)+(in_buffer[16]<<10)+(in_buffer[16]<<11))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<2)-(in_buffer[17]<<4)-(in_buffer[17]<<7)+(in_buffer[17]<<11))+(0-(in_buffer[18]<<0)-(in_buffer[18]<<3)+(in_buffer[18]<<8)+(in_buffer[18]<<11)+(in_buffer[18]<<12))+(0+(in_buffer[19]<<1)+(in_buffer[19]<<2)-(in_buffer[19]<<5)-(in_buffer[19]<<7)-(in_buffer[19]<<9)+(in_buffer[19]<<11)+(in_buffer[19]<<12))-(0+(in_buffer[20]<<2)+(in_buffer[20]<<4)+(in_buffer[20]<<8)+(in_buffer[20]<<11))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<1)+(in_buffer[21]<<4)+(in_buffer[21]<<6))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<4)-(in_buffer[22]<<7)+(in_buffer[22]<<10))-(0+(in_buffer[23]<<0)+(in_buffer[23]<<1)-(in_buffer[23]<<6)+(in_buffer[23]<<10)+(in_buffer[23]<<14))-(0-(in_buffer[24]<<1)-(in_buffer[24]<<3)+(in_buffer[24]<<6)+(in_buffer[24]<<12))+(0-(in_buffer[25]<<0)+(in_buffer[25]<<3)-(in_buffer[25]<<5)+(in_buffer[25]<<7)+(in_buffer[25]<<8)+(in_buffer[25]<<11))-(0+(in_buffer[26]<<0)-(in_buffer[26]<<2)+(in_buffer[26]<<5)+(in_buffer[26]<<7)+(in_buffer[26]<<8)+(in_buffer[26]<<11)+(in_buffer[26]<<12))-(0+(in_buffer[27]<<0)-(in_buffer[27]<<3)-(in_buffer[27]<<5)-(in_buffer[27]<<7)+(in_buffer[27]<<10)+(in_buffer[27]<<11))-(0+(in_buffer[28]<<2)-(in_buffer[28]<<5)+(in_buffer[28]<<10))+(0+(in_buffer[29]<<4)+(in_buffer[29]<<6)+(in_buffer[29]<<10)+(in_buffer[29]<<13))+(0-(in_buffer[30]<<0)+(in_buffer[30]<<2)+(in_buffer[30]<<3)+(in_buffer[30]<<6)+(in_buffer[30]<<8)+(in_buffer[30]<<10)+(in_buffer[30]<<11))-(0-(in_buffer[31]<<0)-(in_buffer[31]<<2)+(in_buffer[31]<<5)+(in_buffer[31]<<11))+(0-(in_buffer[32]<<2)+(in_buffer[32]<<7)+(in_buffer[32]<<9)+(in_buffer[32]<<10))+(0-(in_buffer[33]<<1)+(in_buffer[33]<<6)+(in_buffer[33]<<8)+(in_buffer[33]<<9))-(0-(in_buffer[34]<<0)-(in_buffer[34]<<3)-(in_buffer[34]<<6)-(in_buffer[34]<<9)+(in_buffer[34]<<12)+(in_buffer[34]<<13))-(0+(in_buffer[35]<<1)+(in_buffer[35]<<6)+(in_buffer[35]<<9)+(in_buffer[35]<<10)+(in_buffer[35]<<13))-(0+(in_buffer[36]<<0)+(in_buffer[36]<<3)+(in_buffer[36]<<7)+(in_buffer[36]<<12))-(0+(in_buffer[37]<<3)+(in_buffer[37]<<4)+(in_buffer[37]<<7)+(in_buffer[37]<<9))+(0+(in_buffer[38]<<2)+(in_buffer[38]<<4)+(in_buffer[38]<<8)+(in_buffer[38]<<11))+(0-(in_buffer[39]<<0)+(in_buffer[39]<<2)+(in_buffer[39]<<3)+(in_buffer[39]<<6)+(in_buffer[39]<<8)+(in_buffer[39]<<10)+(in_buffer[39]<<11))+(0+(in_buffer[40]<<1)+(in_buffer[40]<<4)+(in_buffer[40]<<6)+(in_buffer[40]<<10)+(in_buffer[40]<<11))-(0+(in_buffer[41]<<0)+(in_buffer[41]<<2)+(in_buffer[41]<<6)+(in_buffer[41]<<9))-(0-(in_buffer[42]<<0)+(in_buffer[42]<<10)+(in_buffer[42]<<11))+(0+(in_buffer[43]<<0)-(in_buffer[43]<<2)+(in_buffer[43]<<6)-(in_buffer[43]<<8)+(in_buffer[43]<<12))+(0+(in_buffer[44]<<0)+(in_buffer[44]<<1)-(in_buffer[44]<<7)+(in_buffer[44]<<9)+(in_buffer[44]<<10))-(0-(in_buffer[45]<<0)-(in_buffer[45]<<2)-(in_buffer[45]<<4)-(in_buffer[45]<<6)+(in_buffer[45]<<11)+(in_buffer[45]<<12))-(0+(in_buffer[46]<<0)-(in_buffer[46]<<3)-(in_buffer[46]<<5)-(in_buffer[46]<<7)+(in_buffer[46]<<10)+(in_buffer[46]<<11))-(0+(in_buffer[47]<<0)+(in_buffer[47]<<6)+(in_buffer[47]<<7)+(in_buffer[47]<<11))+(0+(in_buffer[48]<<3)+(in_buffer[48]<<7)-(in_buffer[48]<<10)+(in_buffer[48]<<13))+(0+(in_buffer[49]<<1)-(in_buffer[49]<<3)-(in_buffer[49]<<6)+(in_buffer[49]<<9)+(in_buffer[49]<<11))+(0+(in_buffer[50]<<1)+(in_buffer[50]<<3)-(in_buffer[50]<<5)-(in_buffer[50]<<8)+(in_buffer[50]<<12))-(0+(in_buffer[51]<<1)+(in_buffer[51]<<5)-(in_buffer[51]<<8)+(in_buffer[51]<<11))-(0+(in_buffer[52]<<0)+(in_buffer[52]<<3)+(in_buffer[52]<<5)+(in_buffer[52]<<9)+(in_buffer[52]<<10))-(0+(in_buffer[53]<<0)-(in_buffer[53]<<2)-(in_buffer[53]<<5)+(in_buffer[53]<<8)+(in_buffer[53]<<10))+(0+(in_buffer[54]<<1)+(in_buffer[54]<<3)+(in_buffer[54]<<6)+(in_buffer[54]<<8)+(in_buffer[54]<<11)+(in_buffer[54]<<12))+(0-(in_buffer[55]<<1)+(in_buffer[55]<<5)+(in_buffer[55]<<6)+(in_buffer[55]<<9)+(in_buffer[55]<<13))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<6)+(in_buffer[56]<<7)+(in_buffer[56]<<11))+(0-(in_buffer[57]<<4)-(in_buffer[57]<<6)-(in_buffer[57]<<8)+(in_buffer[57]<<12)+(in_buffer[57]<<13))+(0-(in_buffer[58]<<3)+(in_buffer[58]<<8)+(in_buffer[58]<<10)+(in_buffer[58]<<11))+(0+(in_buffer[59]<<0)+(in_buffer[59]<<2)-(in_buffer[59]<<4)-(in_buffer[59]<<7)+(in_buffer[59]<<11))+(0+(in_buffer[60]<<2)+(in_buffer[60]<<4)+(in_buffer[60]<<8)+(in_buffer[60]<<11))+(0-(in_buffer[61]<<0)+(in_buffer[61]<<3)+(in_buffer[61]<<4)+(in_buffer[61]<<7)-(in_buffer[61]<<9)+(in_buffer[61]<<12))-(0+(in_buffer[62]<<0)+(in_buffer[62]<<2)-(in_buffer[62]<<4)-(in_buffer[62]<<7)+(in_buffer[62]<<11))+(0-(in_buffer[63]<<2)-(in_buffer[63]<<4)-(in_buffer[63]<<6)+(in_buffer[63]<<10)+(in_buffer[63]<<11))+(0-(in_buffer[64]<<1)-(in_buffer[64]<<3)-(in_buffer[64]<<5)+(in_buffer[64]<<9)+(in_buffer[64]<<10))+(0-(in_buffer[65]<<3)+(in_buffer[65]<<8)+(in_buffer[65]<<10)+(in_buffer[65]<<11))-(0-(in_buffer[66]<<0)+(in_buffer[66]<<5)+(in_buffer[66]<<7)+(in_buffer[66]<<8))-(0+(in_buffer[67]<<2)+(in_buffer[67]<<4)+(in_buffer[67]<<5)+(in_buffer[67]<<11)+(in_buffer[67]<<13))+(0-(in_buffer[68]<<3)-(in_buffer[68]<<6)+(in_buffer[68]<<9)+(in_buffer[68]<<13))+(0-(in_buffer[69]<<0)+(in_buffer[69]<<3)-(in_buffer[69]<<5)+(in_buffer[69]<<7)+(in_buffer[69]<<8)+(in_buffer[69]<<11))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<1)-(in_buffer[70]<<7)+(in_buffer[70]<<9)+(in_buffer[70]<<10))+(0-(in_buffer[71]<<1)+(in_buffer[71]<<5)-(in_buffer[71]<<7)-(in_buffer[71]<<9)+(in_buffer[71]<<12))+(0-(in_buffer[72]<<2)-(in_buffer[72]<<4)-(in_buffer[72]<<6)+(in_buffer[72]<<10)+(in_buffer[72]<<11))+(0+(in_buffer[73]<<1)+(in_buffer[73]<<2)+(in_buffer[73]<<5)+(in_buffer[73]<<7))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6)-(in_buffer[74]<<8)+(in_buffer[74]<<12))+(0+(in_buffer[75]<<0)-(in_buffer[75]<<2)-(in_buffer[75]<<5)+(in_buffer[75]<<8)+(in_buffer[75]<<10))-(0+(in_buffer[76]<<0)+(in_buffer[76]<<4)-(in_buffer[76]<<7)+(in_buffer[76]<<10))-(0+(in_buffer[77]<<1)+(in_buffer[77]<<3)+(in_buffer[77]<<7)+(in_buffer[77]<<10))-(0+(in_buffer[78]<<0)+(in_buffer[78]<<1)-(in_buffer[78]<<4)-(in_buffer[78]<<7)+(in_buffer[78]<<13))+(0+(in_buffer[79]<<3)+(in_buffer[79]<<5)+(in_buffer[79]<<9)+(in_buffer[79]<<12))-(0-(in_buffer[80]<<1)-(in_buffer[80]<<4)+(in_buffer[80]<<7)+(in_buffer[80]<<11))-(0-(in_buffer[81]<<2)-(in_buffer[81]<<4)-(in_buffer[81]<<6)+(in_buffer[81]<<10)+(in_buffer[81]<<11))-(0+(in_buffer[82]<<4)+(in_buffer[82]<<5)+(in_buffer[82]<<8)+(in_buffer[82]<<10))-(0+(in_buffer[83]<<0)+(in_buffer[83]<<4)-(in_buffer[83]<<7)+(in_buffer[83]<<10))-(0+(in_buffer[84]<<5)+(in_buffer[84]<<6)+(in_buffer[84]<<9)+(in_buffer[84]<<11))+(0-(in_buffer[85]<<0)+(in_buffer[85]<<4)-(in_buffer[85]<<6)-(in_buffer[85]<<8)+(in_buffer[85]<<11))-(0-(in_buffer[86]<<0)+(in_buffer[86]<<3)+(in_buffer[86]<<4)+(in_buffer[86]<<7)-(in_buffer[86]<<9)+(in_buffer[86]<<12))+(0+(in_buffer[87]<<2)+(in_buffer[87]<<3)+(in_buffer[87]<<6)+(in_buffer[87]<<8))+(0-(in_buffer[88]<<1)+(in_buffer[88]<<6)+(in_buffer[88]<<8)+(in_buffer[88]<<9))-(0+(in_buffer[89]<<1)+(in_buffer[89]<<3)+(in_buffer[89]<<7)+(in_buffer[89]<<10))+(0+(in_buffer[90]<<0)+(in_buffer[90]<<1)-(in_buffer[90]<<4)-(in_buffer[90]<<7)+(in_buffer[90]<<13))-(0+(in_buffer[91]<<0)+(in_buffer[91]<<3)+(in_buffer[91]<<5)+(in_buffer[91]<<9)+(in_buffer[91]<<10))-(0+(in_buffer[92]<<0)+(in_buffer[92]<<1)+(in_buffer[92]<<6)+(in_buffer[92]<<9)+(in_buffer[92]<<11)+(in_buffer[92]<<12))-(0+(in_buffer[93]<<1)+(in_buffer[93]<<4)+(in_buffer[93]<<6)+(in_buffer[93]<<10)+(in_buffer[93]<<11))+(0+(in_buffer[94]<<0)+(in_buffer[94]<<6)+(in_buffer[94]<<7)+(in_buffer[94]<<11))-(0+(in_buffer[95]<<0)+(in_buffer[95]<<1)+(in_buffer[95]<<4)+(in_buffer[95]<<6))-(0+(in_buffer[96]<<1)+(in_buffer[96]<<3)+(in_buffer[96]<<7)+(in_buffer[96]<<10))-(0+(in_buffer[97]<<0)-(in_buffer[97]<<2)-(in_buffer[97]<<4)+(in_buffer[97]<<7)+(in_buffer[97]<<10)+(in_buffer[97]<<12))-(0+(in_buffer[98]<<5)+(in_buffer[98]<<6)+(in_buffer[98]<<9)+(in_buffer[98]<<11))+(0+(in_buffer[99]<<2)-(in_buffer[99]<<5)+(in_buffer[99]<<10))-(0+(in_buffer[100]<<0)+(in_buffer[100]<<3)+(in_buffer[100]<<5)+(in_buffer[100]<<9)+(in_buffer[100]<<10))+(0+(in_buffer[101]<<0)+(in_buffer[101]<<2)+(in_buffer[101]<<5)+(in_buffer[101]<<7)+(in_buffer[101]<<10)+(in_buffer[101]<<11))-(0+(in_buffer[102]<<0)-(in_buffer[102]<<2)-(in_buffer[102]<<5)+(in_buffer[102]<<8)+(in_buffer[102]<<10))-(0+(in_buffer[103]<<0)+(in_buffer[103]<<2)+(in_buffer[103]<<5)+(in_buffer[103]<<7)+(in_buffer[103]<<10)+(in_buffer[103]<<11))-(0-(in_buffer[105]<<2)+(in_buffer[105]<<7)+(in_buffer[105]<<9)+(in_buffer[105]<<10))-(0+(in_buffer[106]<<1)-(in_buffer[106]<<4)+(in_buffer[106]<<9))+(0-(in_buffer[107]<<0)+(in_buffer[107]<<3)-(in_buffer[107]<<5)+(in_buffer[107]<<7)+(in_buffer[107]<<8)+(in_buffer[107]<<11))+(0+(in_buffer[108]<<0)+(in_buffer[108]<<4)-(in_buffer[108]<<7)+(in_buffer[108]<<10))+(0+(in_buffer[110]<<0)-(in_buffer[110]<<2)+(in_buffer[110]<<4)+(in_buffer[110]<<5)+(in_buffer[110]<<8)+(in_buffer[110]<<11)+(in_buffer[110]<<13))-(0+(in_buffer[111]<<1)-(in_buffer[111]<<3)-(in_buffer[111]<<6)+(in_buffer[111]<<9)+(in_buffer[111]<<11))+(0+(in_buffer[112]<<0)+(in_buffer[112]<<3)+(in_buffer[112]<<5)+(in_buffer[112]<<9)+(in_buffer[112]<<10))-(0-(in_buffer[113]<<1)-(in_buffer[113]<<4)+(in_buffer[113]<<7)+(in_buffer[113]<<11))-(0-(in_buffer[114]<<0)+(in_buffer[114]<<5)+(in_buffer[114]<<7)+(in_buffer[114]<<8))-(0+(in_buffer[115]<<2)+(in_buffer[115]<<3)+(in_buffer[115]<<6)+(in_buffer[115]<<8))-(0-(in_buffer[116]<<1)+(in_buffer[116]<<11)+(in_buffer[116]<<12))-(0+(in_buffer[117]<<5)-(in_buffer[117]<<8)+(in_buffer[117]<<13))-(0-(in_buffer[118]<<1)-(in_buffer[118]<<3)-(in_buffer[118]<<5)+(in_buffer[118]<<9)+(in_buffer[118]<<10))-(0+(in_buffer[119]<<1)+(in_buffer[119]<<2)+(in_buffer[119]<<5)+(in_buffer[119]<<7))+(0-(in_buffer[120]<<0)+(in_buffer[120]<<3)-(in_buffer[120]<<6)+(in_buffer[120]<<10)+(in_buffer[120]<<12));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight26;
assign in_buffer_weight26=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<7)+(in_buffer[0]<<12))-(0-(in_buffer[1]<<1)-(in_buffer[1]<<3)+(in_buffer[1]<<6)+(in_buffer[1]<<12))-(0+(in_buffer[2]<<0)+(in_buffer[2]<<5)+(in_buffer[2]<<8)+(in_buffer[2]<<9)+(in_buffer[2]<<12))-(0+(in_buffer[3]<<5)+(in_buffer[3]<<6)+(in_buffer[3]<<9)+(in_buffer[3]<<11))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<3)-(in_buffer[4]<<6)-(in_buffer[4]<<8)+(in_buffer[4]<<13))+(0+(in_buffer[5]<<0)-(in_buffer[5]<<3)-(in_buffer[5]<<5)+(in_buffer[5]<<8)+(in_buffer[5]<<10)+(in_buffer[5]<<12)+(in_buffer[5]<<13))+(0-(in_buffer[6]<<3)+(in_buffer[6]<<7)-(in_buffer[6]<<9)-(in_buffer[6]<<11)+(in_buffer[6]<<14))+(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)-(in_buffer[7]<<4)+(in_buffer[7]<<8)+(in_buffer[7]<<9))-(0+(in_buffer[8]<<5)+(in_buffer[8]<<6)+(in_buffer[8]<<9)+(in_buffer[8]<<11))-(0-(in_buffer[9]<<1)-(in_buffer[9]<<4)+(in_buffer[9]<<7)+(in_buffer[9]<<11))+(0+(in_buffer[10]<<2)+(in_buffer[10]<<4)-(in_buffer[10]<<6)-(in_buffer[10]<<9)+(in_buffer[10]<<13))+(0+(in_buffer[11]<<6)+(in_buffer[11]<<7)+(in_buffer[11]<<10)+(in_buffer[11]<<12))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<6)+(in_buffer[12]<<7)+(in_buffer[12]<<11))+(0+(in_buffer[13]<<2)+(in_buffer[13]<<6)-(in_buffer[13]<<9)+(in_buffer[13]<<12))-(0+(in_buffer[14]<<5)+(in_buffer[14]<<6)+(in_buffer[14]<<9)+(in_buffer[14]<<11))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<4)+(in_buffer[15]<<5)+(in_buffer[15]<<8)+(in_buffer[15]<<12))-(0+(in_buffer[16]<<1)-(in_buffer[16]<<4)+(in_buffer[16]<<9))+(0+(in_buffer[17]<<2)-(in_buffer[17]<<5)+(in_buffer[17]<<10))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<7)+(in_buffer[18]<<8)+(in_buffer[18]<<12))-(0+(in_buffer[19]<<0)-(in_buffer[19]<<3)-(in_buffer[19]<<6)-(in_buffer[19]<<9)+(in_buffer[19]<<11)+(in_buffer[19]<<12))-(0-(in_buffer[20]<<0)+(in_buffer[20]<<5)+(in_buffer[20]<<7)+(in_buffer[20]<<8))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<6)+(in_buffer[21]<<9))+(0-(in_buffer[22]<<1)+(in_buffer[22]<<11)+(in_buffer[22]<<12))+(0-(in_buffer[23]<<3)-(in_buffer[23]<<6)+(in_buffer[23]<<9)+(in_buffer[23]<<13))+(0-(in_buffer[24]<<1)-(in_buffer[24]<<4)+(in_buffer[24]<<9)+(in_buffer[24]<<12)+(in_buffer[24]<<13))+(0+(in_buffer[25]<<2)+(in_buffer[25]<<4)-(in_buffer[25]<<6)-(in_buffer[25]<<9)+(in_buffer[25]<<13))+(0+(in_buffer[26]<<2)+(in_buffer[26]<<3)-(in_buffer[26]<<9)+(in_buffer[26]<<11)+(in_buffer[26]<<12))+(0+(in_buffer[27]<<1)-(in_buffer[27]<<3)-(in_buffer[27]<<6)+(in_buffer[27]<<9)+(in_buffer[27]<<11))-(0+(in_buffer[28]<<0)+(in_buffer[28]<<2)+(in_buffer[28]<<6)+(in_buffer[28]<<9))-(0-(in_buffer[29]<<1)-(in_buffer[29]<<4)+(in_buffer[29]<<7)+(in_buffer[29]<<11))-(0+(in_buffer[30]<<1)+(in_buffer[30]<<3)+(in_buffer[30]<<7)+(in_buffer[30]<<10))-(0-(in_buffer[31]<<0)+(in_buffer[31]<<10)+(in_buffer[31]<<11))+(0+(in_buffer[32]<<0)+(in_buffer[32]<<2)+(in_buffer[32]<<6)+(in_buffer[32]<<9))+(0+(in_buffer[33]<<0)-(in_buffer[33]<<3)+(in_buffer[33]<<7)+(in_buffer[33]<<9)+(in_buffer[33]<<11)+(in_buffer[33]<<13))+(0+(in_buffer[34]<<0)+(in_buffer[34]<<2)+(in_buffer[34]<<4)+(in_buffer[34]<<5)-(in_buffer[34]<<10)+(in_buffer[34]<<13))+(0-(in_buffer[35]<<0)-(in_buffer[35]<<2)+(in_buffer[35]<<6)-(in_buffer[35]<<8)+(in_buffer[35]<<11)+(in_buffer[35]<<13))+(0+(in_buffer[36]<<1)-(in_buffer[36]<<5)-(in_buffer[36]<<10)+(in_buffer[36]<<13))+(0+(in_buffer[37]<<0)-(in_buffer[37]<<2)+(in_buffer[37]<<10)+(in_buffer[37]<<13))-(0+(in_buffer[38]<<0)+(in_buffer[38]<<1)-(in_buffer[38]<<4)-(in_buffer[38]<<6)-(in_buffer[38]<<8)+(in_buffer[38]<<10)+(in_buffer[38]<<11))+(0+(in_buffer[39]<<0)+(in_buffer[39]<<2)-(in_buffer[39]<<4)-(in_buffer[39]<<7)+(in_buffer[39]<<11))-(0+(in_buffer[40]<<2)+(in_buffer[40]<<3)+(in_buffer[40]<<6)+(in_buffer[40]<<8))-(0+(in_buffer[41]<<0)+(in_buffer[41]<<1)-(in_buffer[41]<<7)+(in_buffer[41]<<9)+(in_buffer[41]<<10))-(0+(in_buffer[42]<<1)+(in_buffer[42]<<5)-(in_buffer[42]<<8)+(in_buffer[42]<<11))-(0-(in_buffer[43]<<1)+(in_buffer[43]<<6)+(in_buffer[43]<<8)+(in_buffer[43]<<9))+(0+(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<10)+(in_buffer[44]<<13))-(0+(in_buffer[45]<<3)+(in_buffer[45]<<4)+(in_buffer[45]<<7)+(in_buffer[45]<<9))+(0+(in_buffer[46]<<5)+(in_buffer[46]<<6)+(in_buffer[46]<<9)+(in_buffer[46]<<11))+(0-(in_buffer[47]<<0)+(in_buffer[47]<<5)+(in_buffer[47]<<7)+(in_buffer[47]<<8))+(0+(in_buffer[48]<<0)-(in_buffer[48]<<2)-(in_buffer[48]<<4)+(in_buffer[48]<<7)+(in_buffer[48]<<10)+(in_buffer[48]<<12))-(0-(in_buffer[49]<<1)+(in_buffer[49]<<6)+(in_buffer[49]<<8)+(in_buffer[49]<<9))+(0+(in_buffer[50]<<1)+(in_buffer[50]<<5)-(in_buffer[50]<<8)+(in_buffer[50]<<11))+(0+(in_buffer[51]<<0)+(in_buffer[51]<<2)-(in_buffer[51]<<4)-(in_buffer[51]<<7)+(in_buffer[51]<<11))+(0-(in_buffer[52]<<0)+(in_buffer[52]<<5)+(in_buffer[52]<<6)-(in_buffer[52]<<9)+(in_buffer[52]<<11)+(in_buffer[52]<<12))-(0+(in_buffer[54]<<0)+(in_buffer[54]<<3)+(in_buffer[54]<<7)+(in_buffer[54]<<12))-(0-(in_buffer[55]<<0)-(in_buffer[55]<<2)+(in_buffer[55]<<7)+(in_buffer[55]<<9)+(in_buffer[55]<<12))+(0+(in_buffer[56]<<0)+(in_buffer[56]<<3)+(in_buffer[56]<<5)+(in_buffer[56]<<9)+(in_buffer[56]<<10))-(0-(in_buffer[57]<<0)-(in_buffer[57]<<2)-(in_buffer[57]<<4)+(in_buffer[57]<<8)+(in_buffer[57]<<9))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<3)+(in_buffer[58]<<5)+(in_buffer[58]<<9)+(in_buffer[58]<<10))+(0-(in_buffer[59]<<1)-(in_buffer[59]<<3)+(in_buffer[59]<<6)+(in_buffer[59]<<12))-(0-(in_buffer[60]<<0)-(in_buffer[60]<<3)+(in_buffer[60]<<6)+(in_buffer[60]<<10))+(0+(in_buffer[61]<<0)-(in_buffer[61]<<2)+(in_buffer[61]<<6)-(in_buffer[61]<<8)+(in_buffer[61]<<12))-(0+(in_buffer[62]<<0)+(in_buffer[62]<<4)-(in_buffer[62]<<7)+(in_buffer[62]<<10))+(0+(in_buffer[63]<<2)+(in_buffer[63]<<4)+(in_buffer[63]<<8)+(in_buffer[63]<<11))-(0+(in_buffer[64]<<4)-(in_buffer[64]<<7)+(in_buffer[64]<<12))-(0-(in_buffer[65]<<0)+(in_buffer[65]<<5)+(in_buffer[65]<<7)+(in_buffer[65]<<8))-(0-(in_buffer[66]<<3)+(in_buffer[66]<<8)+(in_buffer[66]<<10)+(in_buffer[66]<<11))+(0+(in_buffer[67]<<1)-(in_buffer[67]<<5)-(in_buffer[67]<<10)+(in_buffer[67]<<13))-(0+(in_buffer[68]<<2)+(in_buffer[68]<<3)+(in_buffer[68]<<6)+(in_buffer[68]<<8))-(0-(in_buffer[69]<<1)+(in_buffer[69]<<6)+(in_buffer[69]<<8)+(in_buffer[69]<<9))+(0-(in_buffer[70]<<0)-(in_buffer[70]<<2)+(in_buffer[70]<<7)+(in_buffer[70]<<9)+(in_buffer[70]<<12))-(0+(in_buffer[71]<<1)-(in_buffer[71]<<3)-(in_buffer[71]<<6)+(in_buffer[71]<<9)+(in_buffer[71]<<11))+(0+(in_buffer[72]<<0)+(in_buffer[72]<<6)+(in_buffer[72]<<7)+(in_buffer[72]<<11))-(0-(in_buffer[73]<<1)+(in_buffer[73]<<4)-(in_buffer[73]<<6)+(in_buffer[73]<<8)+(in_buffer[73]<<9)+(in_buffer[73]<<12))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<3)+(in_buffer[74]<<8))+(0+(in_buffer[75]<<0)-(in_buffer[75]<<3)+(in_buffer[75]<<8))+(0-(in_buffer[76]<<0)-(in_buffer[76]<<3)+(in_buffer[76]<<6)+(in_buffer[76]<<10))-(0+(in_buffer[77]<<3)+(in_buffer[77]<<4)+(in_buffer[77]<<7)+(in_buffer[77]<<9))+(0-(in_buffer[78]<<2)+(in_buffer[78]<<7)+(in_buffer[78]<<9)+(in_buffer[78]<<10))-(0+(in_buffer[79]<<2)+(in_buffer[79]<<3)+(in_buffer[79]<<6)+(in_buffer[79]<<8))+(0+(in_buffer[80]<<3)+(in_buffer[80]<<4)+(in_buffer[80]<<7)+(in_buffer[80]<<9))+(0-(in_buffer[81]<<0)-(in_buffer[81]<<2)-(in_buffer[81]<<4)-(in_buffer[81]<<6)+(in_buffer[81]<<11)+(in_buffer[81]<<12))-(0+(in_buffer[82]<<5)+(in_buffer[82]<<6)+(in_buffer[82]<<9)+(in_buffer[82]<<11))+(0+(in_buffer[83]<<0)+(in_buffer[83]<<2)+(in_buffer[83]<<5)+(in_buffer[83]<<7)+(in_buffer[83]<<10)+(in_buffer[83]<<11))-(0+(in_buffer[84]<<4)-(in_buffer[84]<<7)+(in_buffer[84]<<12))+(0+(in_buffer[85]<<0)+(in_buffer[85]<<3)+(in_buffer[85]<<5)+(in_buffer[85]<<9)+(in_buffer[85]<<10))-(0+(in_buffer[86]<<2)+(in_buffer[86]<<3)+(in_buffer[86]<<6)+(in_buffer[86]<<8))-(0+(in_buffer[87]<<1)-(in_buffer[87]<<4)+(in_buffer[87]<<9))+(0+(in_buffer[88]<<1)-(in_buffer[88]<<3)-(in_buffer[88]<<6)+(in_buffer[88]<<9)+(in_buffer[88]<<11))+(0+(in_buffer[89]<<0)-(in_buffer[89]<<4)-(in_buffer[89]<<9)+(in_buffer[89]<<12))+(0-(in_buffer[90]<<1)+(in_buffer[90]<<6)+(in_buffer[90]<<8)+(in_buffer[90]<<9))-(0+(in_buffer[91]<<1)+(in_buffer[91]<<3)-(in_buffer[91]<<5)-(in_buffer[91]<<8)+(in_buffer[91]<<12))+(0-(in_buffer[92]<<0)-(in_buffer[92]<<3)+(in_buffer[92]<<8)+(in_buffer[92]<<11)+(in_buffer[92]<<12))+(0+(in_buffer[93]<<1)+(in_buffer[93]<<2)+(in_buffer[93]<<5)+(in_buffer[93]<<7))+(0+(in_buffer[94]<<1)+(in_buffer[94]<<2)+(in_buffer[94]<<5)+(in_buffer[94]<<7))-(0+(in_buffer[95]<<4)+(in_buffer[95]<<5)+(in_buffer[95]<<8)+(in_buffer[95]<<10))+(0+(in_buffer[96]<<2)+(in_buffer[96]<<4)+(in_buffer[96]<<8)+(in_buffer[96]<<11))+(0+(in_buffer[97]<<1)+(in_buffer[97]<<3)-(in_buffer[97]<<5)-(in_buffer[97]<<8)+(in_buffer[97]<<12))+(0-(in_buffer[98]<<1)+(in_buffer[98]<<5)-(in_buffer[98]<<7)-(in_buffer[98]<<9)+(in_buffer[98]<<12))+(0+(in_buffer[99]<<0)+(in_buffer[99]<<1)-(in_buffer[99]<<5)+(in_buffer[99]<<12))+(0+(in_buffer[100]<<1)+(in_buffer[100]<<4)+(in_buffer[100]<<8)+(in_buffer[100]<<13))+(0-(in_buffer[101]<<2)-(in_buffer[101]<<4)-(in_buffer[101]<<6)+(in_buffer[101]<<10)+(in_buffer[101]<<11))-(0-(in_buffer[102]<<1)+(in_buffer[102]<<3)+(in_buffer[102]<<4)+(in_buffer[102]<<7)+(in_buffer[102]<<9)+(in_buffer[102]<<11)+(in_buffer[102]<<12))+(0-(in_buffer[103]<<2)-(in_buffer[103]<<5)+(in_buffer[103]<<8)+(in_buffer[103]<<12))+(0+(in_buffer[104]<<1)+(in_buffer[104]<<2)+(in_buffer[104]<<5)+(in_buffer[104]<<7))+(0+(in_buffer[105]<<1)+(in_buffer[105]<<2)-(in_buffer[105]<<5)-(in_buffer[105]<<7)-(in_buffer[105]<<9)+(in_buffer[105]<<11)+(in_buffer[105]<<12))-(0+(in_buffer[106]<<0)-(in_buffer[106]<<4)-(in_buffer[106]<<9)+(in_buffer[106]<<12))-(0+(in_buffer[107]<<0)+(in_buffer[107]<<3)+(in_buffer[107]<<7)+(in_buffer[107]<<12))+(0+(in_buffer[108]<<0)+(in_buffer[108]<<1)-(in_buffer[108]<<4)-(in_buffer[108]<<6)-(in_buffer[108]<<8)+(in_buffer[108]<<10)+(in_buffer[108]<<11))-(0+(in_buffer[110]<<0)+(in_buffer[110]<<2)-(in_buffer[110]<<4)-(in_buffer[110]<<7)+(in_buffer[110]<<11))+(0+(in_buffer[111]<<0)+(in_buffer[111]<<4)-(in_buffer[111]<<7)+(in_buffer[111]<<10))+(0+(in_buffer[112]<<0)+(in_buffer[112]<<5)+(in_buffer[112]<<8)+(in_buffer[112]<<9)+(in_buffer[112]<<12))+(0-(in_buffer[113]<<1)-(in_buffer[113]<<3)-(in_buffer[113]<<5)+(in_buffer[113]<<9)+(in_buffer[113]<<10))+(0+(in_buffer[114]<<3)+(in_buffer[114]<<4)+(in_buffer[114]<<7)+(in_buffer[114]<<9))-(0+(in_buffer[115]<<0)+(in_buffer[115]<<1)+(in_buffer[115]<<4)+(in_buffer[115]<<8)+(in_buffer[115]<<10)+(in_buffer[115]<<12))+(0-(in_buffer[116]<<3)-(in_buffer[116]<<6)+(in_buffer[116]<<9)+(in_buffer[116]<<13))+(0+(in_buffer[117]<<1)-(in_buffer[117]<<3)-(in_buffer[117]<<6)+(in_buffer[117]<<9)+(in_buffer[117]<<11))-(0+(in_buffer[118]<<2)+(in_buffer[118]<<3)+(in_buffer[118]<<6)+(in_buffer[118]<<8))+(0+(in_buffer[119]<<1)-(in_buffer[119]<<4)+(in_buffer[119]<<9))-(0-(in_buffer[120]<<0)+(in_buffer[120]<<3)-(in_buffer[120]<<5)+(in_buffer[120]<<7)+(in_buffer[120]<<8)+(in_buffer[120]<<11));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight27;
assign in_buffer_weight27=0+(0-(in_buffer[0]<<1)+(in_buffer[0]<<6)+(in_buffer[0]<<8)+(in_buffer[0]<<9))+(0+(in_buffer[1]<<1)-(in_buffer[1]<<4)+(in_buffer[1]<<9))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<1)+(in_buffer[2]<<4)+(in_buffer[2]<<6))+(0-(in_buffer[3]<<1)+(in_buffer[3]<<6)+(in_buffer[3]<<8)+(in_buffer[3]<<9))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<6)+(in_buffer[4]<<9))+(0-(in_buffer[7]<<0)+(in_buffer[7]<<5)+(in_buffer[7]<<7)+(in_buffer[7]<<8))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<4)-(in_buffer[8]<<7)+(in_buffer[8]<<10))-(0-(in_buffer[9]<<1)+(in_buffer[9]<<6)+(in_buffer[9]<<8)+(in_buffer[9]<<9))-(0+(in_buffer[10]<<1)-(in_buffer[10]<<4)+(in_buffer[10]<<9))-(0+(in_buffer[11]<<0)-(in_buffer[11]<<3)+(in_buffer[11]<<8))+(0+(in_buffer[12]<<1)+(in_buffer[12]<<2)+(in_buffer[12]<<5)+(in_buffer[12]<<7))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<1)+(in_buffer[14]<<4)+(in_buffer[14]<<6))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<1)+(in_buffer[15]<<4)+(in_buffer[15]<<6))+(0-(in_buffer[16]<<0)-(in_buffer[16]<<2)-(in_buffer[16]<<4)+(in_buffer[16]<<8)+(in_buffer[16]<<9))-(0+(in_buffer[17]<<1)-(in_buffer[17]<<4)+(in_buffer[17]<<9))-(0+(in_buffer[18]<<1)+(in_buffer[18]<<2)+(in_buffer[18]<<5)+(in_buffer[18]<<7))+(0+(in_buffer[20]<<3)+(in_buffer[20]<<4)+(in_buffer[20]<<7)+(in_buffer[20]<<9))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<6)+(in_buffer[21]<<9))-(0+(in_buffer[22]<<1)-(in_buffer[22]<<4)+(in_buffer[22]<<9))-(0-(in_buffer[23]<<0)+(in_buffer[23]<<5)+(in_buffer[23]<<7)+(in_buffer[23]<<8))-(0-(in_buffer[24]<<0)+(in_buffer[24]<<5)+(in_buffer[24]<<7)+(in_buffer[24]<<8))-(0-(in_buffer[25]<<0)+(in_buffer[25]<<5)+(in_buffer[25]<<7)+(in_buffer[25]<<8))-(0+(in_buffer[26]<<0)-(in_buffer[26]<<3)+(in_buffer[26]<<8))+(0+(in_buffer[27]<<2)+(in_buffer[27]<<3)+(in_buffer[27]<<6)+(in_buffer[27]<<8))-(0+(in_buffer[28]<<3)+(in_buffer[28]<<4)+(in_buffer[28]<<7)+(in_buffer[28]<<9))+(0-(in_buffer[29]<<0)-(in_buffer[29]<<2)-(in_buffer[29]<<4)+(in_buffer[29]<<8)+(in_buffer[29]<<9))+(0+(in_buffer[30]<<2)+(in_buffer[30]<<3)+(in_buffer[30]<<6)+(in_buffer[30]<<8))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<1)+(in_buffer[31]<<4)+(in_buffer[31]<<6))+(0+(in_buffer[32]<<0)+(in_buffer[32]<<2)+(in_buffer[32]<<6)+(in_buffer[32]<<9))+(0+(in_buffer[33]<<0)-(in_buffer[33]<<3)+(in_buffer[33]<<8))+(0+(in_buffer[34]<<3)+(in_buffer[34]<<4)+(in_buffer[34]<<7)+(in_buffer[34]<<9))-(0+(in_buffer[35]<<2)+(in_buffer[35]<<3)+(in_buffer[35]<<6)+(in_buffer[35]<<8))+(0+(in_buffer[36]<<1)+(in_buffer[36]<<2)+(in_buffer[36]<<5)+(in_buffer[36]<<7))-(0-(in_buffer[37]<<0)+(in_buffer[37]<<5)+(in_buffer[37]<<7)+(in_buffer[37]<<8))-(0+(in_buffer[38]<<0)+(in_buffer[38]<<4)-(in_buffer[38]<<7)+(in_buffer[38]<<10))+(0-(in_buffer[40]<<0)+(in_buffer[40]<<5)+(in_buffer[40]<<7)+(in_buffer[40]<<8))-(0+(in_buffer[41]<<2)+(in_buffer[41]<<3)+(in_buffer[41]<<6)+(in_buffer[41]<<8))+(0+(in_buffer[42]<<3)+(in_buffer[42]<<4)+(in_buffer[42]<<7)+(in_buffer[42]<<9))+(0-(in_buffer[43]<<0)+(in_buffer[43]<<5)+(in_buffer[43]<<7)+(in_buffer[43]<<8))-(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)-(in_buffer[44]<<4)+(in_buffer[44]<<8)+(in_buffer[44]<<9))+(0+(in_buffer[46]<<0)+(in_buffer[46]<<1)+(in_buffer[46]<<4)+(in_buffer[46]<<6))+(0+(in_buffer[47]<<1)+(in_buffer[47]<<2)+(in_buffer[47]<<5)+(in_buffer[47]<<7))+(0+(in_buffer[48]<<0)+(in_buffer[48]<<2)+(in_buffer[48]<<6)+(in_buffer[48]<<9))+(0+(in_buffer[49]<<3)+(in_buffer[49]<<4)+(in_buffer[49]<<7)+(in_buffer[49]<<9))-(0+(in_buffer[50]<<3)+(in_buffer[50]<<4)+(in_buffer[50]<<7)+(in_buffer[50]<<9))+(0+(in_buffer[51]<<1)+(in_buffer[51]<<2)+(in_buffer[51]<<5)+(in_buffer[51]<<7))-(0+(in_buffer[52]<<2)+(in_buffer[52]<<3)+(in_buffer[52]<<6)+(in_buffer[52]<<8))+(0+(in_buffer[53]<<2)+(in_buffer[53]<<3)+(in_buffer[53]<<6)+(in_buffer[53]<<8))-(0+(in_buffer[54]<<3)+(in_buffer[54]<<4)+(in_buffer[54]<<7)+(in_buffer[54]<<9))+(0-(in_buffer[55]<<0)+(in_buffer[55]<<5)+(in_buffer[55]<<7)+(in_buffer[55]<<8))+(0-(in_buffer[56]<<1)+(in_buffer[56]<<6)+(in_buffer[56]<<8)+(in_buffer[56]<<9))-(0-(in_buffer[57]<<1)+(in_buffer[57]<<6)+(in_buffer[57]<<8)+(in_buffer[57]<<9))-(0+(in_buffer[58]<<3)+(in_buffer[58]<<4)+(in_buffer[58]<<7)+(in_buffer[58]<<9))+(0-(in_buffer[59]<<0)+(in_buffer[59]<<5)+(in_buffer[59]<<7)+(in_buffer[59]<<8))+(0+(in_buffer[60]<<0)-(in_buffer[60]<<3)+(in_buffer[60]<<8))+(0-(in_buffer[61]<<1)+(in_buffer[61]<<6)+(in_buffer[61]<<8)+(in_buffer[61]<<9))-(0+(in_buffer[62]<<3)+(in_buffer[62]<<4)+(in_buffer[62]<<7)+(in_buffer[62]<<9))-(0-(in_buffer[63]<<0)-(in_buffer[63]<<2)-(in_buffer[63]<<4)+(in_buffer[63]<<8)+(in_buffer[63]<<9))+(0+(in_buffer[64]<<3)+(in_buffer[64]<<4)+(in_buffer[64]<<7)+(in_buffer[64]<<9))+(0-(in_buffer[67]<<0)-(in_buffer[67]<<2)-(in_buffer[67]<<4)+(in_buffer[67]<<8)+(in_buffer[67]<<9))-(0+(in_buffer[68]<<0)-(in_buffer[68]<<3)+(in_buffer[68]<<8))-(0+(in_buffer[70]<<0)+(in_buffer[70]<<4)-(in_buffer[70]<<7)+(in_buffer[70]<<10))-(0+(in_buffer[71]<<0)+(in_buffer[71]<<2)+(in_buffer[71]<<6)+(in_buffer[71]<<9))-(0+(in_buffer[72]<<2)+(in_buffer[72]<<3)+(in_buffer[72]<<6)+(in_buffer[72]<<8))+(0+(in_buffer[73]<<2)+(in_buffer[73]<<3)+(in_buffer[73]<<6)+(in_buffer[73]<<8))-(0+(in_buffer[74]<<2)+(in_buffer[74]<<3)+(in_buffer[74]<<6)+(in_buffer[74]<<8))-(0+(in_buffer[75]<<2)+(in_buffer[75]<<3)+(in_buffer[75]<<6)+(in_buffer[75]<<8))+(0+(in_buffer[76]<<3)+(in_buffer[76]<<4)+(in_buffer[76]<<7)+(in_buffer[76]<<9))+(0-(in_buffer[77]<<0)+(in_buffer[77]<<5)+(in_buffer[77]<<7)+(in_buffer[77]<<8))-(0+(in_buffer[78]<<1)+(in_buffer[78]<<2)+(in_buffer[78]<<5)+(in_buffer[78]<<7))-(0+(in_buffer[79]<<1)+(in_buffer[79]<<2)+(in_buffer[79]<<5)+(in_buffer[79]<<7))-(0+(in_buffer[80]<<2)+(in_buffer[80]<<3)+(in_buffer[80]<<6)+(in_buffer[80]<<8))-(0+(in_buffer[81]<<3)+(in_buffer[81]<<4)+(in_buffer[81]<<7)+(in_buffer[81]<<9))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)-(in_buffer[82]<<4)+(in_buffer[82]<<8)+(in_buffer[82]<<9))+(0-(in_buffer[83]<<1)+(in_buffer[83]<<6)+(in_buffer[83]<<8)+(in_buffer[83]<<9))-(0-(in_buffer[84]<<0)+(in_buffer[84]<<5)+(in_buffer[84]<<7)+(in_buffer[84]<<8))+(0+(in_buffer[86]<<2)+(in_buffer[86]<<3)+(in_buffer[86]<<6)+(in_buffer[86]<<8))-(0-(in_buffer[87]<<0)-(in_buffer[87]<<2)-(in_buffer[87]<<4)+(in_buffer[87]<<8)+(in_buffer[87]<<9))-(0+(in_buffer[88]<<1)+(in_buffer[88]<<2)+(in_buffer[88]<<5)+(in_buffer[88]<<7))-(0+(in_buffer[89]<<1)+(in_buffer[89]<<2)+(in_buffer[89]<<5)+(in_buffer[89]<<7))+(0+(in_buffer[90]<<0)+(in_buffer[90]<<2)+(in_buffer[90]<<6)+(in_buffer[90]<<9))-(0+(in_buffer[91]<<3)+(in_buffer[91]<<4)+(in_buffer[91]<<7)+(in_buffer[91]<<9))-(0+(in_buffer[92]<<2)+(in_buffer[92]<<3)+(in_buffer[92]<<6)+(in_buffer[92]<<8))+(0+(in_buffer[93]<<0)+(in_buffer[93]<<1)+(in_buffer[93]<<4)+(in_buffer[93]<<6))-(0+(in_buffer[95]<<0)+(in_buffer[95]<<1)+(in_buffer[95]<<4)+(in_buffer[95]<<6))-(0+(in_buffer[96]<<0)+(in_buffer[96]<<4)-(in_buffer[96]<<7)+(in_buffer[96]<<10))+(0+(in_buffer[97]<<1)+(in_buffer[97]<<2)+(in_buffer[97]<<5)+(in_buffer[97]<<7))+(0-(in_buffer[98]<<0)-(in_buffer[98]<<2)-(in_buffer[98]<<4)+(in_buffer[98]<<8)+(in_buffer[98]<<9))-(0+(in_buffer[99]<<2)+(in_buffer[99]<<3)+(in_buffer[99]<<6)+(in_buffer[99]<<8))-(0+(in_buffer[100]<<3)+(in_buffer[100]<<4)+(in_buffer[100]<<7)+(in_buffer[100]<<9))-(0+(in_buffer[101]<<0)-(in_buffer[101]<<3)+(in_buffer[101]<<8))-(0+(in_buffer[102]<<0)+(in_buffer[102]<<4)-(in_buffer[102]<<7)+(in_buffer[102]<<10))-(0+(in_buffer[104]<<0)+(in_buffer[104]<<1)+(in_buffer[104]<<4)+(in_buffer[104]<<6))-(0+(in_buffer[105]<<1)-(in_buffer[105]<<4)+(in_buffer[105]<<9))-(0+(in_buffer[106]<<0)+(in_buffer[106]<<2)+(in_buffer[106]<<6)+(in_buffer[106]<<9))-(0+(in_buffer[108]<<0)+(in_buffer[108]<<1)+(in_buffer[108]<<4)+(in_buffer[108]<<6))-(0+(in_buffer[109]<<0)+(in_buffer[109]<<1)+(in_buffer[109]<<4)+(in_buffer[109]<<6))-(0+(in_buffer[112]<<1)+(in_buffer[112]<<2)+(in_buffer[112]<<5)+(in_buffer[112]<<7))-(0+(in_buffer[114]<<0)+(in_buffer[114]<<1)+(in_buffer[114]<<4)+(in_buffer[114]<<6))-(0+(in_buffer[115]<<2)+(in_buffer[115]<<3)+(in_buffer[115]<<6)+(in_buffer[115]<<8))+(0-(in_buffer[117]<<1)+(in_buffer[117]<<6)+(in_buffer[117]<<8)+(in_buffer[117]<<9))-(0+(in_buffer[118]<<3)+(in_buffer[118]<<4)+(in_buffer[118]<<7)+(in_buffer[118]<<9))-(0+(in_buffer[119]<<0)-(in_buffer[119]<<3)+(in_buffer[119]<<8))+(0+(in_buffer[120]<<0)+(in_buffer[120]<<4)-(in_buffer[120]<<7)+(in_buffer[120]<<10));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight28;
assign in_buffer_weight28=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<3)+(in_buffer[0]<<7)+(in_buffer[0]<<12))+(0-(in_buffer[1]<<0)+(in_buffer[1]<<5)+(in_buffer[1]<<6)-(in_buffer[1]<<9)+(in_buffer[1]<<11)+(in_buffer[1]<<12))-(0+(in_buffer[2]<<0)-(in_buffer[2]<<3)-(in_buffer[2]<<5)-(in_buffer[2]<<7)+(in_buffer[2]<<10)+(in_buffer[2]<<11))-(0+(in_buffer[3]<<1)+(in_buffer[3]<<2)-(in_buffer[3]<<5)-(in_buffer[3]<<8)+(in_buffer[3]<<14))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<1)-(in_buffer[4]<<7)+(in_buffer[4]<<9)+(in_buffer[4]<<10))+(0+(in_buffer[5]<<6)-(in_buffer[5]<<9)+(in_buffer[5]<<14))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<5)+(in_buffer[6]<<7)+(in_buffer[6]<<10)+(in_buffer[6]<<11))-(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)+(in_buffer[7]<<4)+(in_buffer[7]<<5)+(in_buffer[7]<<8)+(in_buffer[7]<<14))-(0+(in_buffer[8]<<6)+(in_buffer[8]<<7)+(in_buffer[8]<<10)+(in_buffer[8]<<12))+(0+(in_buffer[9]<<3)-(in_buffer[9]<<6)+(in_buffer[9]<<11))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)-(in_buffer[10]<<4)-(in_buffer[10]<<7)+(in_buffer[10]<<13))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<4)+(in_buffer[11]<<6)+(in_buffer[11]<<11)+(in_buffer[11]<<12))-(0+(in_buffer[12]<<0)+(in_buffer[12]<<5)+(in_buffer[12]<<8)+(in_buffer[12]<<9)+(in_buffer[12]<<12))+(0-(in_buffer[13]<<0)+(in_buffer[13]<<5)+(in_buffer[13]<<7)+(in_buffer[13]<<8))+(0-(in_buffer[14]<<1)+(in_buffer[14]<<5)-(in_buffer[14]<<7)-(in_buffer[14]<<9)+(in_buffer[14]<<12))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<4)-(in_buffer[15]<<7)+(in_buffer[15]<<10))+(0-(in_buffer[16]<<2)-(in_buffer[16]<<4)+(in_buffer[16]<<7)+(in_buffer[16]<<13))+(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)-(in_buffer[17]<<4)+(in_buffer[17]<<8)+(in_buffer[17]<<9))+(0+(in_buffer[18]<<1)-(in_buffer[18]<<4)+(in_buffer[18]<<9))+(0+(in_buffer[19]<<1)-(in_buffer[19]<<3)-(in_buffer[19]<<6)+(in_buffer[19]<<9)+(in_buffer[19]<<11))-(0-(in_buffer[20]<<0)-(in_buffer[20]<<2)-(in_buffer[20]<<5)+(in_buffer[20]<<8)-(in_buffer[20]<<10)+(in_buffer[20]<<13))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<1)+(in_buffer[21]<<6)+(in_buffer[21]<<9)+(in_buffer[21]<<11)+(in_buffer[21]<<12))-(0+(in_buffer[22]<<2)-(in_buffer[22]<<4)-(in_buffer[22]<<7)+(in_buffer[22]<<10)+(in_buffer[22]<<12))-(0+(in_buffer[23]<<1)-(in_buffer[23]<<4)-(in_buffer[23]<<6)-(in_buffer[23]<<8)+(in_buffer[23]<<11)+(in_buffer[23]<<12))-(0+(in_buffer[25]<<0)+(in_buffer[25]<<3)+(in_buffer[25]<<5)+(in_buffer[25]<<9)+(in_buffer[25]<<10))-(0+(in_buffer[26]<<5)+(in_buffer[26]<<6)+(in_buffer[26]<<9)+(in_buffer[26]<<11))+(0+(in_buffer[27]<<0)-(in_buffer[27]<<4)-(in_buffer[27]<<9)+(in_buffer[27]<<12))-(0-(in_buffer[28]<<0)+(in_buffer[28]<<3)-(in_buffer[28]<<5)+(in_buffer[28]<<7)+(in_buffer[28]<<8)+(in_buffer[28]<<11))-(0-(in_buffer[29]<<0)+(in_buffer[29]<<5)+(in_buffer[29]<<6)-(in_buffer[29]<<9)+(in_buffer[29]<<11)+(in_buffer[29]<<12))+(0+(in_buffer[30]<<0)+(in_buffer[30]<<1)-(in_buffer[30]<<4)-(in_buffer[30]<<6)-(in_buffer[30]<<8)+(in_buffer[30]<<10)+(in_buffer[30]<<11))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<2)-(in_buffer[31]<<8)+(in_buffer[31]<<11)+(in_buffer[31]<<12))+(0+(in_buffer[32]<<2)+(in_buffer[32]<<3)+(in_buffer[32]<<6)+(in_buffer[32]<<8))-(0-(in_buffer[33]<<1)-(in_buffer[33]<<4)-(in_buffer[33]<<7)-(in_buffer[33]<<10)+(in_buffer[33]<<13)+(in_buffer[33]<<14))-(0+(in_buffer[34]<<1)+(in_buffer[34]<<5)-(in_buffer[34]<<8)+(in_buffer[34]<<11))+(0+(in_buffer[35]<<2)-(in_buffer[35]<<5)+(in_buffer[35]<<10))+(0-(in_buffer[36]<<1)+(in_buffer[36]<<6)+(in_buffer[36]<<8)+(in_buffer[36]<<9))-(0-(in_buffer[37]<<3)-(in_buffer[37]<<5)-(in_buffer[37]<<7)+(in_buffer[37]<<11)+(in_buffer[37]<<12))+(0-(in_buffer[38]<<0)+(in_buffer[38]<<3)-(in_buffer[38]<<6)+(in_buffer[38]<<10)+(in_buffer[38]<<12))-(0+(in_buffer[39]<<3)+(in_buffer[39]<<4)+(in_buffer[39]<<7)+(in_buffer[39]<<9))-(0+(in_buffer[40]<<1)-(in_buffer[40]<<4)+(in_buffer[40]<<9))+(0+(in_buffer[41]<<6)+(in_buffer[41]<<7)+(in_buffer[41]<<10)+(in_buffer[41]<<12))-(0-(in_buffer[42]<<0)+(in_buffer[42]<<3)+(in_buffer[42]<<4)+(in_buffer[42]<<7)-(in_buffer[42]<<9)+(in_buffer[42]<<12))+(0+(in_buffer[43]<<0)+(in_buffer[43]<<1)-(in_buffer[43]<<7)+(in_buffer[43]<<9)+(in_buffer[43]<<10))-(0-(in_buffer[44]<<1)+(in_buffer[44]<<6)-(in_buffer[44]<<9)-(in_buffer[44]<<11)+(in_buffer[44]<<13)+(in_buffer[44]<<14))-(0-(in_buffer[45]<<3)-(in_buffer[45]<<5)-(in_buffer[45]<<7)+(in_buffer[45]<<11)+(in_buffer[45]<<12))-(0+(in_buffer[46]<<0)+(in_buffer[46]<<3)+(in_buffer[46]<<5)+(in_buffer[46]<<9)+(in_buffer[46]<<10))-(0+(in_buffer[47]<<0)+(in_buffer[47]<<2)+(in_buffer[47]<<6)+(in_buffer[47]<<9))-(0+(in_buffer[48]<<4)+(in_buffer[48]<<6)+(in_buffer[48]<<10)+(in_buffer[48]<<13))+(0+(in_buffer[49]<<0)+(in_buffer[49]<<1)-(in_buffer[49]<<7)+(in_buffer[49]<<9)+(in_buffer[49]<<10))+(0+(in_buffer[50]<<3)+(in_buffer[50]<<4)+(in_buffer[50]<<7)+(in_buffer[50]<<9))+(0+(in_buffer[51]<<0)-(in_buffer[51]<<4)-(in_buffer[51]<<9)+(in_buffer[51]<<12))+(0+(in_buffer[52]<<0)-(in_buffer[52]<<2)-(in_buffer[52]<<4)+(in_buffer[52]<<7)+(in_buffer[52]<<10)+(in_buffer[52]<<12))+(0+(in_buffer[53]<<3)-(in_buffer[53]<<6)+(in_buffer[53]<<11))+(0+(in_buffer[54]<<1)-(in_buffer[54]<<3)-(in_buffer[54]<<6)+(in_buffer[54]<<9)+(in_buffer[54]<<11))-(0-(in_buffer[55]<<1)-(in_buffer[55]<<3)+(in_buffer[55]<<6)+(in_buffer[55]<<12))-(0-(in_buffer[56]<<0)-(in_buffer[56]<<3)-(in_buffer[56]<<5)-(in_buffer[56]<<7)+(in_buffer[56]<<10)+(in_buffer[56]<<13))+(0+(in_buffer[58]<<0)+(in_buffer[58]<<1)-(in_buffer[58]<<7)+(in_buffer[58]<<9)+(in_buffer[58]<<10))-(0+(in_buffer[59]<<0)+(in_buffer[59]<<1)-(in_buffer[59]<<7)+(in_buffer[59]<<9)+(in_buffer[59]<<10))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)-(in_buffer[60]<<7)+(in_buffer[60]<<9)+(in_buffer[60]<<10))-(0+(in_buffer[61]<<0)+(in_buffer[61]<<5)+(in_buffer[61]<<8)+(in_buffer[61]<<9)+(in_buffer[61]<<12))+(0-(in_buffer[62]<<0)+(in_buffer[62]<<4)-(in_buffer[62]<<6)-(in_buffer[62]<<8)+(in_buffer[62]<<11))+(0+(in_buffer[63]<<2)+(in_buffer[63]<<4)+(in_buffer[63]<<8)+(in_buffer[63]<<11))-(0+(in_buffer[64]<<3)-(in_buffer[64]<<6)+(in_buffer[64]<<11))-(0+(in_buffer[65]<<1)+(in_buffer[65]<<2)-(in_buffer[65]<<5)-(in_buffer[65]<<7)-(in_buffer[65]<<9)+(in_buffer[65]<<11)+(in_buffer[65]<<12))-(0+(in_buffer[66]<<1)+(in_buffer[66]<<4)+(in_buffer[66]<<6)+(in_buffer[66]<<10)+(in_buffer[66]<<11))-(0-(in_buffer[67]<<0)+(in_buffer[67]<<5)+(in_buffer[67]<<7)+(in_buffer[67]<<8))+(0+(in_buffer[68]<<5)+(in_buffer[68]<<6)+(in_buffer[68]<<9)+(in_buffer[68]<<11))+(0+(in_buffer[69]<<1)-(in_buffer[69]<<4)+(in_buffer[69]<<9))-(0+(in_buffer[70]<<0)+(in_buffer[70]<<6)+(in_buffer[70]<<7)+(in_buffer[70]<<11))+(0+(in_buffer[71]<<1)+(in_buffer[71]<<2)+(in_buffer[71]<<5)+(in_buffer[71]<<7))-(0+(in_buffer[72]<<0)+(in_buffer[72]<<1)-(in_buffer[72]<<7)+(in_buffer[72]<<9)+(in_buffer[72]<<10))+(0+(in_buffer[73]<<1)+(in_buffer[73]<<4)+(in_buffer[73]<<6)+(in_buffer[73]<<10)+(in_buffer[73]<<11))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<4)-(in_buffer[74]<<9)+(in_buffer[74]<<12))-(0+(in_buffer[75]<<1)+(in_buffer[75]<<3)+(in_buffer[75]<<7)+(in_buffer[75]<<10))-(0-(in_buffer[76]<<0)+(in_buffer[76]<<10)+(in_buffer[76]<<11))-(0+(in_buffer[77]<<0)+(in_buffer[77]<<2)+(in_buffer[77]<<6)+(in_buffer[77]<<9))+(0+(in_buffer[78]<<5)-(in_buffer[78]<<8)+(in_buffer[78]<<13))+(0+(in_buffer[79]<<0)+(in_buffer[79]<<1)-(in_buffer[79]<<4)-(in_buffer[79]<<6)-(in_buffer[79]<<8)+(in_buffer[79]<<10)+(in_buffer[79]<<11))+(0-(in_buffer[80]<<0)+(in_buffer[80]<<5)+(in_buffer[80]<<7)+(in_buffer[80]<<8))+(0+(in_buffer[81]<<1)+(in_buffer[81]<<3)+(in_buffer[81]<<7)+(in_buffer[81]<<10))+(0-(in_buffer[82]<<0)-(in_buffer[82]<<2)+(in_buffer[82]<<5)+(in_buffer[82]<<11))+(0+(in_buffer[83]<<0)+(in_buffer[83]<<4)-(in_buffer[83]<<7)+(in_buffer[83]<<10))-(0+(in_buffer[84]<<0)+(in_buffer[84]<<3)+(in_buffer[84]<<5)+(in_buffer[84]<<9)+(in_buffer[84]<<10))+(0+(in_buffer[85]<<0)+(in_buffer[85]<<4)-(in_buffer[85]<<7)+(in_buffer[85]<<10))+(0+(in_buffer[86]<<1)+(in_buffer[86]<<3)+(in_buffer[86]<<6)+(in_buffer[86]<<8)+(in_buffer[86]<<11)+(in_buffer[86]<<12))-(0+(in_buffer[87]<<1)+(in_buffer[87]<<5)-(in_buffer[87]<<8)+(in_buffer[87]<<11))-(0+(in_buffer[88]<<0)+(in_buffer[88]<<2)+(in_buffer[88]<<4)+(in_buffer[88]<<5)-(in_buffer[88]<<10)+(in_buffer[88]<<13))+(0+(in_buffer[89]<<1)+(in_buffer[89]<<7)+(in_buffer[89]<<8)+(in_buffer[89]<<12))+(0+(in_buffer[90]<<0)-(in_buffer[90]<<2)-(in_buffer[90]<<5)+(in_buffer[90]<<8)+(in_buffer[90]<<10))+(0+(in_buffer[91]<<1)+(in_buffer[91]<<3)+(in_buffer[91]<<7)+(in_buffer[91]<<10))+(0+(in_buffer[92]<<0)+(in_buffer[92]<<2)+(in_buffer[92]<<3)+(in_buffer[92]<<9)+(in_buffer[92]<<11))+(0+(in_buffer[93]<<0)-(in_buffer[93]<<3)+(in_buffer[93]<<8))-(0-(in_buffer[94]<<0)-(in_buffer[94]<<2)+(in_buffer[94]<<7)+(in_buffer[94]<<9)+(in_buffer[94]<<12))-(0-(in_buffer[95]<<1)+(in_buffer[95]<<11)+(in_buffer[95]<<12))+(0+(in_buffer[96]<<1)+(in_buffer[96]<<3)+(in_buffer[96]<<7)+(in_buffer[96]<<10))+(0+(in_buffer[97]<<0)-(in_buffer[97]<<2)+(in_buffer[97]<<10)+(in_buffer[97]<<13))+(0+(in_buffer[98]<<0)+(in_buffer[98]<<2)+(in_buffer[98]<<6)+(in_buffer[98]<<9))-(0+(in_buffer[99]<<2)-(in_buffer[99]<<4)-(in_buffer[99]<<7)+(in_buffer[99]<<10)+(in_buffer[99]<<12))+(0-(in_buffer[100]<<1)+(in_buffer[100]<<5)-(in_buffer[100]<<7)-(in_buffer[100]<<9)+(in_buffer[100]<<12))-(0+(in_buffer[101]<<0)+(in_buffer[101]<<2)+(in_buffer[101]<<3)+(in_buffer[101]<<9)+(in_buffer[101]<<11))+(0-(in_buffer[102]<<1)+(in_buffer[102]<<4)-(in_buffer[102]<<6)+(in_buffer[102]<<8)+(in_buffer[102]<<9)+(in_buffer[102]<<12))+(0+(in_buffer[103]<<2)+(in_buffer[103]<<4)+(in_buffer[103]<<8)+(in_buffer[103]<<11))+(0+(in_buffer[104]<<0)+(in_buffer[104]<<6)+(in_buffer[104]<<7)+(in_buffer[104]<<11))-(0-(in_buffer[105]<<1)+(in_buffer[105]<<5)-(in_buffer[105]<<7)-(in_buffer[105]<<9)+(in_buffer[105]<<12))-(0+(in_buffer[106]<<0)+(in_buffer[106]<<2)+(in_buffer[106]<<6)+(in_buffer[106]<<9))-(0+(in_buffer[107]<<5)+(in_buffer[107]<<6)+(in_buffer[107]<<9)+(in_buffer[107]<<11))+(0-(in_buffer[108]<<1)+(in_buffer[108]<<4)+(in_buffer[108]<<5)+(in_buffer[108]<<8)-(in_buffer[108]<<10)+(in_buffer[108]<<13))+(0+(in_buffer[109]<<1)+(in_buffer[109]<<4)+(in_buffer[109]<<6)+(in_buffer[109]<<10)+(in_buffer[109]<<11))-(0+(in_buffer[110]<<6)+(in_buffer[110]<<7)+(in_buffer[110]<<10)+(in_buffer[110]<<12))+(0-(in_buffer[111]<<0)-(in_buffer[111]<<2)-(in_buffer[111]<<4)+(in_buffer[111]<<7)-(in_buffer[111]<<10)+(in_buffer[111]<<12)+(in_buffer[111]<<13))-(0-(in_buffer[112]<<0)-(in_buffer[112]<<2)-(in_buffer[112]<<4)-(in_buffer[112]<<6)+(in_buffer[112]<<11)+(in_buffer[112]<<12))-(0+(in_buffer[113]<<2)-(in_buffer[113]<<6)-(in_buffer[113]<<11)+(in_buffer[113]<<14))+(0-(in_buffer[114]<<2)-(in_buffer[114]<<4)-(in_buffer[114]<<6)+(in_buffer[114]<<10)+(in_buffer[114]<<11))+(0+(in_buffer[115]<<0)-(in_buffer[115]<<3)-(in_buffer[115]<<5)-(in_buffer[115]<<7)+(in_buffer[115]<<10)+(in_buffer[115]<<11))+(0-(in_buffer[116]<<0)+(in_buffer[116]<<10)+(in_buffer[116]<<11))-(0+(in_buffer[117]<<1)+(in_buffer[117]<<3)+(in_buffer[117]<<5)-(in_buffer[117]<<7)+(in_buffer[117]<<10)+(in_buffer[117]<<13))-(0+(in_buffer[118]<<2)+(in_buffer[118]<<4)+(in_buffer[118]<<5)+(in_buffer[118]<<11)+(in_buffer[118]<<13))+(0+(in_buffer[119]<<1)+(in_buffer[119]<<2)+(in_buffer[119]<<7)+(in_buffer[119]<<10)+(in_buffer[119]<<12)+(in_buffer[119]<<13))+(0+(in_buffer[120]<<3)+(in_buffer[120]<<4)+(in_buffer[120]<<7)+(in_buffer[120]<<9));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight29;
assign in_buffer_weight29=0-(0-(in_buffer[0]<<1)-(in_buffer[0]<<4)-(in_buffer[0]<<6)-(in_buffer[0]<<8)+(in_buffer[0]<<11)+(in_buffer[0]<<14))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<3)+(in_buffer[1]<<5)+(in_buffer[1]<<6)+(in_buffer[1]<<10)+(in_buffer[1]<<14))-(0+(in_buffer[2]<<0)+(in_buffer[2]<<2)+(in_buffer[2]<<3)+(in_buffer[2]<<9)+(in_buffer[2]<<11))+(0+(in_buffer[3]<<2)+(in_buffer[3]<<4)+(in_buffer[3]<<8)+(in_buffer[3]<<11))+(0+(in_buffer[4]<<0)-(in_buffer[4]<<2)+(in_buffer[4]<<5)+(in_buffer[4]<<7)+(in_buffer[4]<<8)+(in_buffer[4]<<11)+(in_buffer[4]<<12))+(0+(in_buffer[5]<<1)+(in_buffer[5]<<2)+(in_buffer[5]<<5)+(in_buffer[5]<<7))+(0+(in_buffer[6]<<3)+(in_buffer[6]<<5)+(in_buffer[6]<<9)+(in_buffer[6]<<12))+(0+(in_buffer[7]<<0)-(in_buffer[7]<<3)-(in_buffer[7]<<5)-(in_buffer[7]<<7)+(in_buffer[7]<<10)+(in_buffer[7]<<11))-(0+(in_buffer[8]<<6)+(in_buffer[8]<<7)+(in_buffer[8]<<10)+(in_buffer[8]<<12))-(0+(in_buffer[9]<<0)-(in_buffer[9]<<3)+(in_buffer[9]<<10)+(in_buffer[9]<<12)+(in_buffer[9]<<14))-(0-(in_buffer[10]<<0)+(in_buffer[10]<<3)-(in_buffer[10]<<7)-(in_buffer[10]<<10)+(in_buffer[10]<<15))-(0-(in_buffer[11]<<0)+(in_buffer[11]<<3)+(in_buffer[11]<<5)+(in_buffer[11]<<8)-(in_buffer[11]<<12)+(in_buffer[11]<<15))-(0+(in_buffer[12]<<2)+(in_buffer[12]<<4)+(in_buffer[12]<<8)+(in_buffer[12]<<11))-(0-(in_buffer[13]<<0)-(in_buffer[13]<<3)+(in_buffer[13]<<6)+(in_buffer[13]<<10))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<5)+(in_buffer[14]<<7)+(in_buffer[14]<<10)+(in_buffer[14]<<11))+(0+(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<6)+(in_buffer[15]<<9))-(0-(in_buffer[16]<<0)-(in_buffer[16]<<2)-(in_buffer[16]<<4)+(in_buffer[16]<<8)+(in_buffer[16]<<9))-(0-(in_buffer[17]<<0)-(in_buffer[17]<<2)+(in_buffer[17]<<5)+(in_buffer[17]<<11))-(0-(in_buffer[18]<<2)-(in_buffer[18]<<5)+(in_buffer[18]<<8)+(in_buffer[18]<<12))-(0-(in_buffer[19]<<2)-(in_buffer[19]<<5)+(in_buffer[19]<<8)+(in_buffer[19]<<12))-(0+(in_buffer[20]<<7)+(in_buffer[20]<<8)+(in_buffer[20]<<11)+(in_buffer[20]<<13))-(0-(in_buffer[21]<<5)-(in_buffer[21]<<8)+(in_buffer[21]<<11)+(in_buffer[21]<<15))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<2)-(in_buffer[22]<<4)+(in_buffer[22]<<10)+(in_buffer[22]<<15))+(0-(in_buffer[23]<<1)-(in_buffer[23]<<3)+(in_buffer[23]<<6)+(in_buffer[23]<<12))+(0+(in_buffer[24]<<5)-(in_buffer[24]<<8)+(in_buffer[24]<<13))+(0+(in_buffer[25]<<0)+(in_buffer[25]<<2)-(in_buffer[25]<<8)+(in_buffer[25]<<11)+(in_buffer[25]<<12))-(0+(in_buffer[26]<<1)-(in_buffer[26]<<3)-(in_buffer[26]<<6)+(in_buffer[26]<<9)+(in_buffer[26]<<11))-(0+(in_buffer[27]<<0)-(in_buffer[27]<<3)+(in_buffer[27]<<8))+(0+(in_buffer[28]<<0)-(in_buffer[28]<<3)+(in_buffer[28]<<8))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<2)+(in_buffer[29]<<3)-(in_buffer[29]<<6)-(in_buffer[29]<<8)+(in_buffer[29]<<13))-(0-(in_buffer[30]<<2)-(in_buffer[30]<<5)+(in_buffer[30]<<8)+(in_buffer[30]<<12))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<1)-(in_buffer[31]<<6)+(in_buffer[31]<<10)+(in_buffer[31]<<14))-(0+(in_buffer[32]<<0)-(in_buffer[32]<<2)+(in_buffer[32]<<6)+(in_buffer[32]<<7)-(in_buffer[32]<<11)+(in_buffer[32]<<14))-(0-(in_buffer[33]<<1)-(in_buffer[33]<<4)+(in_buffer[33]<<9)+(in_buffer[33]<<12)+(in_buffer[33]<<13))+(0+(in_buffer[34]<<5)+(in_buffer[34]<<6)+(in_buffer[34]<<9)+(in_buffer[34]<<11))+(0+(in_buffer[35]<<1)-(in_buffer[35]<<3)-(in_buffer[35]<<6)+(in_buffer[35]<<9)+(in_buffer[35]<<11))+(0+(in_buffer[36]<<5)+(in_buffer[36]<<6)+(in_buffer[36]<<9)+(in_buffer[36]<<11))-(0+(in_buffer[37]<<1)+(in_buffer[37]<<2)-(in_buffer[37]<<8)+(in_buffer[37]<<10)+(in_buffer[37]<<11))-(0-(in_buffer[38]<<1)+(in_buffer[38]<<11)+(in_buffer[38]<<12))+(0+(in_buffer[39]<<0)+(in_buffer[39]<<2)+(in_buffer[39]<<4)-(in_buffer[39]<<6)+(in_buffer[39]<<9)+(in_buffer[39]<<12))+(0-(in_buffer[40]<<0)+(in_buffer[40]<<4)-(in_buffer[40]<<7)-(in_buffer[40]<<10)+(in_buffer[40]<<13))-(0-(in_buffer[41]<<0)+(in_buffer[41]<<6)+(in_buffer[41]<<7)+(in_buffer[41]<<13))-(0+(in_buffer[42]<<3)-(in_buffer[42]<<6)+(in_buffer[42]<<11))-(0+(in_buffer[43]<<0)+(in_buffer[43]<<2)-(in_buffer[43]<<8)+(in_buffer[43]<<11)+(in_buffer[43]<<12))-(0+(in_buffer[44]<<3)+(in_buffer[44]<<5)+(in_buffer[44]<<9)+(in_buffer[44]<<12))+(0+(in_buffer[45]<<2)+(in_buffer[45]<<4)+(in_buffer[45]<<8)+(in_buffer[45]<<11))-(0+(in_buffer[46]<<0)-(in_buffer[46]<<4)-(in_buffer[46]<<9)+(in_buffer[46]<<12))+(0-(in_buffer[47]<<0)-(in_buffer[47]<<2)+(in_buffer[47]<<7)+(in_buffer[47]<<9)+(in_buffer[47]<<12))+(0+(in_buffer[48]<<0)+(in_buffer[48]<<1)-(in_buffer[48]<<5)+(in_buffer[48]<<12))-(0+(in_buffer[49]<<0)+(in_buffer[49]<<1)-(in_buffer[49]<<7)+(in_buffer[49]<<9)+(in_buffer[49]<<10))+(0-(in_buffer[50]<<2)-(in_buffer[50]<<5)+(in_buffer[50]<<8)+(in_buffer[50]<<12))+(0+(in_buffer[51]<<1)+(in_buffer[51]<<3)+(in_buffer[51]<<7)+(in_buffer[51]<<10))-(0+(in_buffer[52]<<2)+(in_buffer[52]<<5)+(in_buffer[52]<<7)+(in_buffer[52]<<11)+(in_buffer[52]<<12))-(0-(in_buffer[53]<<1)+(in_buffer[53]<<6)+(in_buffer[53]<<8)+(in_buffer[53]<<9))-(0-(in_buffer[54]<<1)-(in_buffer[54]<<4)+(in_buffer[54]<<7)+(in_buffer[54]<<11))-(0+(in_buffer[55]<<2)+(in_buffer[55]<<5)+(in_buffer[55]<<7)+(in_buffer[55]<<11)+(in_buffer[55]<<12))+(0-(in_buffer[56]<<2)+(in_buffer[56]<<7)+(in_buffer[56]<<9)+(in_buffer[56]<<10))-(0-(in_buffer[57]<<0)-(in_buffer[57]<<2)-(in_buffer[57]<<4)+(in_buffer[57]<<8)+(in_buffer[57]<<9))+(0-(in_buffer[58]<<3)+(in_buffer[58]<<8)+(in_buffer[58]<<10)+(in_buffer[58]<<11))-(0-(in_buffer[59]<<1)-(in_buffer[59]<<4)+(in_buffer[59]<<7)+(in_buffer[59]<<11))+(0+(in_buffer[60]<<0)-(in_buffer[60]<<3)+(in_buffer[60]<<8))+(0+(in_buffer[61]<<0)+(in_buffer[61]<<1)-(in_buffer[61]<<7)+(in_buffer[61]<<9)+(in_buffer[61]<<10))-(0-(in_buffer[62]<<0)+(in_buffer[62]<<4)-(in_buffer[62]<<6)-(in_buffer[62]<<8)+(in_buffer[62]<<11))+(0+(in_buffer[64]<<1)+(in_buffer[64]<<5)-(in_buffer[64]<<8)+(in_buffer[64]<<11))+(0+(in_buffer[65]<<1)-(in_buffer[65]<<3)-(in_buffer[65]<<6)+(in_buffer[65]<<9)+(in_buffer[65]<<11))+(0-(in_buffer[66]<<0)+(in_buffer[66]<<3)+(in_buffer[66]<<4)+(in_buffer[66]<<7)-(in_buffer[66]<<9)+(in_buffer[66]<<12))-(0+(in_buffer[67]<<0)+(in_buffer[67]<<2)+(in_buffer[67]<<5)+(in_buffer[67]<<7)+(in_buffer[67]<<10)+(in_buffer[67]<<11))-(0+(in_buffer[68]<<0)+(in_buffer[68]<<6)+(in_buffer[68]<<7)+(in_buffer[68]<<11))+(0-(in_buffer[69]<<0)+(in_buffer[69]<<10)+(in_buffer[69]<<11))+(0+(in_buffer[70]<<0)+(in_buffer[70]<<1)-(in_buffer[70]<<4)-(in_buffer[70]<<6)-(in_buffer[70]<<8)+(in_buffer[70]<<10)+(in_buffer[70]<<11))-(0-(in_buffer[71]<<0)+(in_buffer[71]<<3)-(in_buffer[71]<<5)+(in_buffer[71]<<7)+(in_buffer[71]<<8)+(in_buffer[71]<<11))+(0+(in_buffer[72]<<2)+(in_buffer[72]<<6)-(in_buffer[72]<<9)+(in_buffer[72]<<12))-(0-(in_buffer[73]<<0)+(in_buffer[73]<<4)-(in_buffer[73]<<6)-(in_buffer[73]<<8)+(in_buffer[73]<<11))-(0+(in_buffer[74]<<0)-(in_buffer[74]<<3)+(in_buffer[74]<<8))+(0+(in_buffer[75]<<1)+(in_buffer[75]<<4)+(in_buffer[75]<<6)+(in_buffer[75]<<10)+(in_buffer[75]<<11))-(0+(in_buffer[76]<<3)-(in_buffer[76]<<6)+(in_buffer[76]<<11))+(0-(in_buffer[77]<<0)+(in_buffer[77]<<3)-(in_buffer[77]<<5)+(in_buffer[77]<<7)+(in_buffer[77]<<8)+(in_buffer[77]<<11))-(0-(in_buffer[78]<<1)-(in_buffer[78]<<4)+(in_buffer[78]<<7)+(in_buffer[78]<<11))+(0+(in_buffer[79]<<2)-(in_buffer[79]<<5)+(in_buffer[79]<<10))+(0-(in_buffer[80]<<0)-(in_buffer[80]<<3)+(in_buffer[80]<<6)+(in_buffer[80]<<10))-(0-(in_buffer[81]<<1)+(in_buffer[81]<<6)+(in_buffer[81]<<8)+(in_buffer[81]<<9))-(0+(in_buffer[82]<<0)+(in_buffer[82]<<2)+(in_buffer[82]<<4)-(in_buffer[82]<<6)+(in_buffer[82]<<9)+(in_buffer[82]<<12))+(0+(in_buffer[83]<<1)-(in_buffer[83]<<3)-(in_buffer[83]<<6)+(in_buffer[83]<<9)+(in_buffer[83]<<11))-(0-(in_buffer[84]<<0)-(in_buffer[84]<<2)-(in_buffer[84]<<4)+(in_buffer[84]<<8)+(in_buffer[84]<<9))-(0+(in_buffer[86]<<5)+(in_buffer[86]<<6)+(in_buffer[86]<<9)+(in_buffer[86]<<11))+(0+(in_buffer[87]<<5)+(in_buffer[87]<<6)+(in_buffer[87]<<9)+(in_buffer[87]<<11))-(0+(in_buffer[88]<<0)+(in_buffer[88]<<2)+(in_buffer[88]<<4)+(in_buffer[88]<<5)-(in_buffer[88]<<10)+(in_buffer[88]<<13))-(0+(in_buffer[89]<<6)+(in_buffer[89]<<7)+(in_buffer[89]<<10)+(in_buffer[89]<<12))+(0+(in_buffer[90]<<1)-(in_buffer[90]<<3)-(in_buffer[90]<<6)+(in_buffer[90]<<9)+(in_buffer[90]<<11))-(0-(in_buffer[91]<<0)-(in_buffer[91]<<2)+(in_buffer[91]<<5)+(in_buffer[91]<<11))-(0+(in_buffer[92]<<0)+(in_buffer[92]<<6)+(in_buffer[92]<<7)+(in_buffer[92]<<11))-(0-(in_buffer[93]<<2)+(in_buffer[93]<<7)+(in_buffer[93]<<9)+(in_buffer[93]<<10))+(0-(in_buffer[94]<<0)+(in_buffer[94]<<4)+(in_buffer[94]<<6)+(in_buffer[94]<<12)+(in_buffer[94]<<13))+(0+(in_buffer[95]<<0)-(in_buffer[95]<<7)-(in_buffer[95]<<9)+(in_buffer[95]<<13))+(0-(in_buffer[96]<<1)+(in_buffer[96]<<6)+(in_buffer[96]<<8)+(in_buffer[96]<<9))-(0+(in_buffer[97]<<0)+(in_buffer[97]<<1)-(in_buffer[97]<<4)-(in_buffer[97]<<6)-(in_buffer[97]<<8)+(in_buffer[97]<<10)+(in_buffer[97]<<11))+(0+(in_buffer[98]<<2)+(in_buffer[98]<<4)+(in_buffer[98]<<8)+(in_buffer[98]<<11))-(0-(in_buffer[99]<<0)-(in_buffer[99]<<2)+(in_buffer[99]<<4)+(in_buffer[99]<<5)+(in_buffer[99]<<8)+(in_buffer[99]<<14))-(0-(in_buffer[100]<<0)+(in_buffer[100]<<4)+(in_buffer[100]<<5)+(in_buffer[100]<<8)+(in_buffer[100]<<12))+(0+(in_buffer[101]<<0)+(in_buffer[101]<<1)-(in_buffer[101]<<5)+(in_buffer[101]<<12))-(0-(in_buffer[102]<<1)+(in_buffer[102]<<5)-(in_buffer[102]<<7)-(in_buffer[102]<<9)+(in_buffer[102]<<12))+(0+(in_buffer[103]<<2)-(in_buffer[103]<<5)+(in_buffer[103]<<10))-(0+(in_buffer[104]<<0)+(in_buffer[104]<<1)-(in_buffer[104]<<4)-(in_buffer[104]<<6)-(in_buffer[104]<<8)+(in_buffer[104]<<10)+(in_buffer[104]<<11))+(0-(in_buffer[105]<<1)+(in_buffer[105]<<4)+(in_buffer[105]<<5)+(in_buffer[105]<<8)-(in_buffer[105]<<10)+(in_buffer[105]<<13))+(0+(in_buffer[106]<<0)+(in_buffer[106]<<3)+(in_buffer[106]<<5)+(in_buffer[106]<<9)+(in_buffer[106]<<10))+(0-(in_buffer[107]<<0)-(in_buffer[107]<<3)+(in_buffer[107]<<6)+(in_buffer[107]<<10))-(0-(in_buffer[108]<<2)-(in_buffer[108]<<4)-(in_buffer[108]<<6)+(in_buffer[108]<<10)+(in_buffer[108]<<11))-(0+(in_buffer[109]<<3)+(in_buffer[109]<<9)+(in_buffer[109]<<10)+(in_buffer[109]<<14))-(0+(in_buffer[110]<<1)+(in_buffer[110]<<3)-(in_buffer[110]<<9)+(in_buffer[110]<<12)+(in_buffer[110]<<13))+(0+(in_buffer[111]<<2)+(in_buffer[111]<<3)-(in_buffer[111]<<9)+(in_buffer[111]<<11)+(in_buffer[111]<<12))+(0+(in_buffer[112]<<5)+(in_buffer[112]<<6)+(in_buffer[112]<<9)+(in_buffer[112]<<11))-(0-(in_buffer[113]<<1)+(in_buffer[113]<<6)+(in_buffer[113]<<7)-(in_buffer[113]<<10)+(in_buffer[113]<<12)+(in_buffer[113]<<13))-(0+(in_buffer[114]<<1)+(in_buffer[114]<<2)-(in_buffer[114]<<5)-(in_buffer[114]<<7)-(in_buffer[114]<<9)+(in_buffer[114]<<11)+(in_buffer[114]<<12))-(0+(in_buffer[115]<<0)-(in_buffer[115]<<3)+(in_buffer[115]<<7)+(in_buffer[115]<<9)+(in_buffer[115]<<11)+(in_buffer[115]<<13))+(0+(in_buffer[116]<<1)+(in_buffer[116]<<3)+(in_buffer[116]<<7)+(in_buffer[116]<<10))-(0+(in_buffer[117]<<0)+(in_buffer[117]<<2)+(in_buffer[117]<<3)+(in_buffer[117]<<9)+(in_buffer[117]<<11))+(0+(in_buffer[118]<<0)-(in_buffer[118]<<2)+(in_buffer[118]<<6)-(in_buffer[118]<<8)+(in_buffer[118]<<12))+(0-(in_buffer[119]<<0)+(in_buffer[119]<<5)-(in_buffer[119]<<8)-(in_buffer[119]<<10)+(in_buffer[119]<<12)+(in_buffer[119]<<13))-(0-(in_buffer[120]<<0)-(in_buffer[120]<<2)-(in_buffer[120]<<4)+(in_buffer[120]<<7)-(in_buffer[120]<<10)+(in_buffer[120]<<12)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight30;
assign in_buffer_weight30=0-(0-(in_buffer[0]<<0)-(in_buffer[0]<<2)-(in_buffer[0]<<4)+(in_buffer[0]<<8)+(in_buffer[0]<<9))+(0+(in_buffer[1]<<3)+(in_buffer[1]<<6)+(in_buffer[1]<<8)+(in_buffer[1]<<12)+(in_buffer[1]<<13))-(0+(in_buffer[2]<<3)+(in_buffer[2]<<5)+(in_buffer[2]<<9)+(in_buffer[2]<<12))-(0-(in_buffer[3]<<2)-(in_buffer[3]<<4)-(in_buffer[3]<<6)+(in_buffer[3]<<10)+(in_buffer[3]<<11))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)-(in_buffer[4]<<4)-(in_buffer[4]<<7)+(in_buffer[4]<<11))+(0+(in_buffer[5]<<0)-(in_buffer[5]<<3)-(in_buffer[5]<<5)-(in_buffer[5]<<7)+(in_buffer[5]<<10)+(in_buffer[5]<<11))-(0+(in_buffer[6]<<0)-(in_buffer[6]<<3)-(in_buffer[6]<<5)-(in_buffer[6]<<7)+(in_buffer[6]<<10)+(in_buffer[6]<<11))-(0+(in_buffer[7]<<1)+(in_buffer[7]<<3)+(in_buffer[7]<<7)+(in_buffer[7]<<10))+(0+(in_buffer[8]<<4)+(in_buffer[8]<<5)+(in_buffer[8]<<8)+(in_buffer[8]<<10))+(0+(in_buffer[9]<<0)-(in_buffer[9]<<3)+(in_buffer[9]<<6)-(in_buffer[9]<<8)+(in_buffer[9]<<14))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)+(in_buffer[10]<<4)+(in_buffer[10]<<8)+(in_buffer[10]<<10)+(in_buffer[10]<<12))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<4)+(in_buffer[11]<<5)-(in_buffer[11]<<10)+(in_buffer[11]<<13))-(0+(in_buffer[12]<<3)+(in_buffer[12]<<9)+(in_buffer[12]<<10)+(in_buffer[12]<<14))-(0+(in_buffer[13]<<1)-(in_buffer[13]<<4)-(in_buffer[13]<<6)-(in_buffer[13]<<8)+(in_buffer[13]<<11)+(in_buffer[13]<<12))+(0+(in_buffer[14]<<0)-(in_buffer[14]<<2)+(in_buffer[14]<<6)-(in_buffer[14]<<8)+(in_buffer[14]<<12))-(0-(in_buffer[15]<<1)-(in_buffer[15]<<3)+(in_buffer[15]<<6)+(in_buffer[15]<<12))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<2)-(in_buffer[16]<<4)-(in_buffer[16]<<7)+(in_buffer[16]<<11))-(0+(in_buffer[17]<<2)+(in_buffer[17]<<4)+(in_buffer[17]<<8)+(in_buffer[17]<<11))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<2)+(in_buffer[18]<<3)+(in_buffer[18]<<9)+(in_buffer[18]<<11))-(0-(in_buffer[19]<<0)+(in_buffer[19]<<4)-(in_buffer[19]<<7)-(in_buffer[19]<<10)+(in_buffer[19]<<13))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<3)-(in_buffer[20]<<5)-(in_buffer[20]<<7)+(in_buffer[20]<<10)+(in_buffer[20]<<11))+(0+(in_buffer[21]<<2)+(in_buffer[21]<<5)+(in_buffer[21]<<7)+(in_buffer[21]<<11)+(in_buffer[21]<<12))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<2)+(in_buffer[22]<<5)-(in_buffer[22]<<9)-(in_buffer[22]<<11)+(in_buffer[22]<<14))-(0-(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<9)+(in_buffer[23]<<13)+(in_buffer[23]<<15))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<1)-(in_buffer[24]<<5)+(in_buffer[24]<<12))+(0+(in_buffer[25]<<2)-(in_buffer[25]<<5)+(in_buffer[25]<<10))-(0+(in_buffer[26]<<0)+(in_buffer[26]<<2)+(in_buffer[26]<<6)+(in_buffer[26]<<9))+(0+(in_buffer[27]<<1)+(in_buffer[27]<<3)+(in_buffer[27]<<7)+(in_buffer[27]<<10))+(0+(in_buffer[28]<<3)+(in_buffer[28]<<4)+(in_buffer[28]<<7)+(in_buffer[28]<<9))+(0+(in_buffer[29]<<0)-(in_buffer[29]<<3)-(in_buffer[29]<<6)-(in_buffer[29]<<9)+(in_buffer[29]<<11)+(in_buffer[29]<<12))-(0+(in_buffer[30]<<3)+(in_buffer[30]<<4)+(in_buffer[30]<<7)+(in_buffer[30]<<9))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<3)+(in_buffer[31]<<4)+(in_buffer[31]<<13))+(0+(in_buffer[32]<<3)+(in_buffer[32]<<5)+(in_buffer[32]<<9)+(in_buffer[32]<<12))-(0+(in_buffer[33]<<0)+(in_buffer[33]<<1)+(in_buffer[33]<<4)+(in_buffer[33]<<6)+(in_buffer[33]<<8)+(in_buffer[33]<<9)+(in_buffer[33]<<12)+(in_buffer[33]<<14))-(0-(in_buffer[34]<<0)-(in_buffer[34]<<3)+(in_buffer[34]<<6)+(in_buffer[34]<<9)+(in_buffer[34]<<11)+(in_buffer[34]<<13)+(in_buffer[34]<<15))+(0-(in_buffer[35]<<0)-(in_buffer[35]<<2)+(in_buffer[35]<<6)-(in_buffer[35]<<8)+(in_buffer[35]<<11)+(in_buffer[35]<<13))-(0+(in_buffer[36]<<2)+(in_buffer[36]<<4)+(in_buffer[36]<<8)+(in_buffer[36]<<11))-(0+(in_buffer[37]<<2)-(in_buffer[37]<<4)-(in_buffer[37]<<7)+(in_buffer[37]<<10)+(in_buffer[37]<<12))-(0+(in_buffer[38]<<1)+(in_buffer[38]<<2)-(in_buffer[38]<<8)+(in_buffer[38]<<10)+(in_buffer[38]<<11))+(0+(in_buffer[40]<<2)+(in_buffer[40]<<6)-(in_buffer[40]<<9)+(in_buffer[40]<<12))+(0-(in_buffer[41]<<0)+(in_buffer[41]<<4)-(in_buffer[41]<<6)-(in_buffer[41]<<8)+(in_buffer[41]<<11))-(0+(in_buffer[42]<<0)+(in_buffer[42]<<4)-(in_buffer[42]<<7)+(in_buffer[42]<<10))+(0-(in_buffer[43]<<0)+(in_buffer[43]<<4)+(in_buffer[43]<<5)+(in_buffer[43]<<8)+(in_buffer[43]<<12))-(0+(in_buffer[44]<<0)+(in_buffer[44]<<2)+(in_buffer[44]<<5)-(in_buffer[44]<<7)+(in_buffer[44]<<13)+(in_buffer[44]<<14))-(0+(in_buffer[45]<<1)-(in_buffer[45]<<3)+(in_buffer[45]<<6)+(in_buffer[45]<<9)+(in_buffer[45]<<10)+(in_buffer[45]<<15))+(0+(in_buffer[46]<<3)+(in_buffer[46]<<7)-(in_buffer[46]<<10)+(in_buffer[46]<<13))-(0+(in_buffer[47]<<5)+(in_buffer[47]<<6)+(in_buffer[47]<<9)+(in_buffer[47]<<11))-(0-(in_buffer[48]<<2)+(in_buffer[48]<<7)+(in_buffer[48]<<9)+(in_buffer[48]<<10))+(0+(in_buffer[49]<<0)-(in_buffer[49]<<2)-(in_buffer[49]<<5)+(in_buffer[49]<<8)+(in_buffer[49]<<10))-(0+(in_buffer[50]<<0)-(in_buffer[50]<<2)-(in_buffer[50]<<5)+(in_buffer[50]<<8)+(in_buffer[50]<<10))+(0-(in_buffer[51]<<1)-(in_buffer[51]<<3)-(in_buffer[51]<<5)+(in_buffer[51]<<9)+(in_buffer[51]<<10))+(0+(in_buffer[52]<<1)-(in_buffer[52]<<5)-(in_buffer[52]<<10)+(in_buffer[52]<<13))-(0+(in_buffer[53]<<2)+(in_buffer[53]<<3)+(in_buffer[53]<<6)+(in_buffer[53]<<8))+(0-(in_buffer[54]<<1)-(in_buffer[54]<<3)+(in_buffer[54]<<8)+(in_buffer[54]<<10)+(in_buffer[54]<<13))-(0+(in_buffer[55]<<2)+(in_buffer[55]<<3)-(in_buffer[55]<<9)+(in_buffer[55]<<11)+(in_buffer[55]<<12))-(0+(in_buffer[56]<<1)+(in_buffer[56]<<2)-(in_buffer[56]<<5)-(in_buffer[56]<<8)+(in_buffer[56]<<14))+(0-(in_buffer[57]<<0)+(in_buffer[57]<<4)-(in_buffer[57]<<6)-(in_buffer[57]<<8)+(in_buffer[57]<<11))-(0+(in_buffer[58]<<2)+(in_buffer[58]<<3)+(in_buffer[58]<<6)+(in_buffer[58]<<8))-(0+(in_buffer[59]<<0)-(in_buffer[59]<<2)-(in_buffer[59]<<5)+(in_buffer[59]<<8)+(in_buffer[59]<<10))+(0-(in_buffer[60]<<0)+(in_buffer[60]<<10)+(in_buffer[60]<<11))+(0-(in_buffer[61]<<0)+(in_buffer[61]<<4)-(in_buffer[61]<<6)-(in_buffer[61]<<8)+(in_buffer[61]<<11))+(0+(in_buffer[62]<<0)+(in_buffer[62]<<2)+(in_buffer[62]<<5)+(in_buffer[62]<<7)+(in_buffer[62]<<10)+(in_buffer[62]<<11))+(0+(in_buffer[63]<<0)-(in_buffer[63]<<4)-(in_buffer[63]<<6)+(in_buffer[63]<<8)+(in_buffer[63]<<9)+(in_buffer[63]<<13))-(0-(in_buffer[64]<<3)+(in_buffer[64]<<8)+(in_buffer[64]<<10)+(in_buffer[64]<<11))+(0+(in_buffer[65]<<0)-(in_buffer[65]<<7)-(in_buffer[65]<<9)+(in_buffer[65]<<13))+(0+(in_buffer[66]<<1)+(in_buffer[66]<<2)-(in_buffer[66]<<6)+(in_buffer[66]<<13))-(0+(in_buffer[67]<<0)+(in_buffer[67]<<1)-(in_buffer[67]<<5)+(in_buffer[67]<<12))-(0-(in_buffer[68]<<2)-(in_buffer[68]<<5)+(in_buffer[68]<<8)+(in_buffer[68]<<12))-(0+(in_buffer[69]<<0)-(in_buffer[69]<<3)-(in_buffer[69]<<5)-(in_buffer[69]<<7)+(in_buffer[69]<<10)+(in_buffer[69]<<11))-(0+(in_buffer[70]<<0)+(in_buffer[70]<<1)-(in_buffer[70]<<7)+(in_buffer[70]<<9)+(in_buffer[70]<<10))+(0+(in_buffer[71]<<1)-(in_buffer[71]<<4)+(in_buffer[71]<<9))+(0-(in_buffer[72]<<0)-(in_buffer[72]<<2)+(in_buffer[72]<<5)+(in_buffer[72]<<11))+(0-(in_buffer[73]<<1)+(in_buffer[73]<<6)+(in_buffer[73]<<8)+(in_buffer[73]<<9))+(0+(in_buffer[74]<<0)-(in_buffer[74]<<2)+(in_buffer[74]<<6)-(in_buffer[74]<<8)+(in_buffer[74]<<12))-(0-(in_buffer[75]<<0)+(in_buffer[75]<<5)+(in_buffer[75]<<6)-(in_buffer[75]<<9)+(in_buffer[75]<<11)+(in_buffer[75]<<12))-(0+(in_buffer[76]<<1)+(in_buffer[76]<<2)+(in_buffer[76]<<5)+(in_buffer[76]<<7))+(0-(in_buffer[77]<<1)+(in_buffer[77]<<4)-(in_buffer[77]<<6)+(in_buffer[77]<<8)+(in_buffer[77]<<9)+(in_buffer[77]<<12))+(0+(in_buffer[78]<<2)-(in_buffer[78]<<5)+(in_buffer[78]<<10))+(0+(in_buffer[79]<<0)+(in_buffer[79]<<1)-(in_buffer[79]<<4)-(in_buffer[79]<<6)-(in_buffer[79]<<8)+(in_buffer[79]<<10)+(in_buffer[79]<<11))-(0-(in_buffer[80]<<0)+(in_buffer[80]<<5)+(in_buffer[80]<<6)-(in_buffer[80]<<9)+(in_buffer[80]<<11)+(in_buffer[80]<<12))+(0+(in_buffer[81]<<0)-(in_buffer[81]<<2)-(in_buffer[81]<<5)+(in_buffer[81]<<8)+(in_buffer[81]<<10))-(0+(in_buffer[82]<<0)-(in_buffer[82]<<3)+(in_buffer[82]<<8))+(0+(in_buffer[83]<<5)+(in_buffer[83]<<6)+(in_buffer[83]<<9)+(in_buffer[83]<<11))-(0-(in_buffer[84]<<2)-(in_buffer[84]<<4)-(in_buffer[84]<<6)+(in_buffer[84]<<10)+(in_buffer[84]<<11))+(0-(in_buffer[85]<<3)+(in_buffer[85]<<8)+(in_buffer[85]<<10)+(in_buffer[85]<<11))-(0-(in_buffer[86]<<2)+(in_buffer[86]<<7)+(in_buffer[86]<<9)+(in_buffer[86]<<10))+(0+(in_buffer[87]<<0)+(in_buffer[87]<<6)+(in_buffer[87]<<7)+(in_buffer[87]<<11))+(0+(in_buffer[88]<<0)-(in_buffer[88]<<2)+(in_buffer[88]<<10)+(in_buffer[88]<<13))+(0+(in_buffer[89]<<0)+(in_buffer[89]<<1)-(in_buffer[89]<<5)+(in_buffer[89]<<12))-(0+(in_buffer[90]<<2)+(in_buffer[90]<<6)-(in_buffer[90]<<9)+(in_buffer[90]<<12))-(0+(in_buffer[91]<<1)+(in_buffer[91]<<2)+(in_buffer[91]<<7)+(in_buffer[91]<<10)+(in_buffer[91]<<12)+(in_buffer[91]<<13))+(0-(in_buffer[92]<<0)-(in_buffer[92]<<2)+(in_buffer[92]<<5)+(in_buffer[92]<<11))+(0+(in_buffer[93]<<0)+(in_buffer[93]<<2)+(in_buffer[93]<<6)+(in_buffer[93]<<9))+(0+(in_buffer[94]<<0)+(in_buffer[94]<<1)+(in_buffer[94]<<6)+(in_buffer[94]<<9)+(in_buffer[94]<<11)+(in_buffer[94]<<12))-(0+(in_buffer[95]<<0)+(in_buffer[95]<<2)-(in_buffer[95]<<8)+(in_buffer[95]<<11)+(in_buffer[95]<<12))-(0+(in_buffer[96]<<0)+(in_buffer[96]<<1)-(in_buffer[96]<<5)+(in_buffer[96]<<12))+(0+(in_buffer[97]<<0)+(in_buffer[97]<<2)-(in_buffer[97]<<8)+(in_buffer[97]<<11)+(in_buffer[97]<<12))+(0-(in_buffer[98]<<0)+(in_buffer[98]<<2)+(in_buffer[98]<<3)+(in_buffer[98]<<9)+(in_buffer[98]<<13))+(0-(in_buffer[99]<<0)+(in_buffer[99]<<6)+(in_buffer[99]<<7)+(in_buffer[99]<<13))-(0-(in_buffer[100]<<3)+(in_buffer[100]<<8)+(in_buffer[100]<<10)+(in_buffer[100]<<11))-(0+(in_buffer[101]<<0)-(in_buffer[101]<<2)-(in_buffer[101]<<4)-(in_buffer[101]<<9)+(in_buffer[101]<<14))-(0+(in_buffer[102]<<0)+(in_buffer[102]<<3)+(in_buffer[102]<<4)+(in_buffer[102]<<13))+(0-(in_buffer[103]<<0)-(in_buffer[103]<<2)-(in_buffer[103]<<5)+(in_buffer[103]<<8)-(in_buffer[103]<<10)+(in_buffer[103]<<13))+(0+(in_buffer[104]<<0)+(in_buffer[104]<<2)-(in_buffer[104]<<8)+(in_buffer[104]<<11)+(in_buffer[104]<<12))+(0+(in_buffer[105]<<1)+(in_buffer[105]<<2)-(in_buffer[105]<<5)-(in_buffer[105]<<7)-(in_buffer[105]<<9)+(in_buffer[105]<<11)+(in_buffer[105]<<12))-(0+(in_buffer[106]<<0)+(in_buffer[106]<<3)+(in_buffer[106]<<7)+(in_buffer[106]<<12))-(0+(in_buffer[107]<<1)-(in_buffer[107]<<3)+(in_buffer[107]<<6)+(in_buffer[107]<<8)+(in_buffer[107]<<9)+(in_buffer[107]<<12)+(in_buffer[107]<<13))-(0+(in_buffer[108]<<0)+(in_buffer[108]<<2)+(in_buffer[108]<<4)-(in_buffer[108]<<6)+(in_buffer[108]<<9)+(in_buffer[108]<<12))+(0-(in_buffer[109]<<1)+(in_buffer[109]<<4)-(in_buffer[109]<<6)+(in_buffer[109]<<8)+(in_buffer[109]<<9)+(in_buffer[109]<<12))-(0+(in_buffer[110]<<0)+(in_buffer[110]<<1)+(in_buffer[110]<<4)+(in_buffer[110]<<6))-(0+(in_buffer[111]<<1)+(in_buffer[111]<<3)+(in_buffer[111]<<5)-(in_buffer[111]<<7)+(in_buffer[111]<<10)+(in_buffer[111]<<13))-(0-(in_buffer[112]<<1)+(in_buffer[112]<<4)+(in_buffer[112]<<6)-(in_buffer[112]<<10)+(in_buffer[112]<<14))+(0+(in_buffer[113]<<1)+(in_buffer[113]<<3)+(in_buffer[113]<<7)+(in_buffer[113]<<10))+(0+(in_buffer[114]<<0)+(in_buffer[114]<<2)+(in_buffer[114]<<3)-(in_buffer[114]<<6)-(in_buffer[114]<<8)+(in_buffer[114]<<13))+(0+(in_buffer[115]<<1)+(in_buffer[115]<<2)+(in_buffer[115]<<5)+(in_buffer[115]<<7))+(0-(in_buffer[116]<<0)-(in_buffer[116]<<2)-(in_buffer[116]<<4)-(in_buffer[116]<<6)+(in_buffer[116]<<11)+(in_buffer[116]<<12))-(0+(in_buffer[117]<<1)+(in_buffer[117]<<2)-(in_buffer[117]<<8)+(in_buffer[117]<<10)+(in_buffer[117]<<11))-(0+(in_buffer[118]<<0)+(in_buffer[118]<<2)-(in_buffer[118]<<8)+(in_buffer[118]<<11)+(in_buffer[118]<<12))-(0+(in_buffer[119]<<0)+(in_buffer[119]<<5)+(in_buffer[119]<<7)-(in_buffer[119]<<10)+(in_buffer[119]<<14))+(0+(in_buffer[120]<<0)-(in_buffer[120]<<7)-(in_buffer[120]<<9)+(in_buffer[120]<<13));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight31;
assign in_buffer_weight31=0-(0+(in_buffer[0]<<3)+(in_buffer[0]<<7)-(in_buffer[0]<<10)+(in_buffer[0]<<13))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)-(in_buffer[1]<<6)-(in_buffer[1]<<10)+(in_buffer[1]<<12)+(in_buffer[1]<<13))-(0+(in_buffer[2]<<1)+(in_buffer[2]<<5)+(in_buffer[2]<<7)+(in_buffer[2]<<12)+(in_buffer[2]<<13))+(0-(in_buffer[3]<<0)+(in_buffer[3]<<3)+(in_buffer[3]<<5)-(in_buffer[3]<<9)+(in_buffer[3]<<13))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<5)+(in_buffer[4]<<7)+(in_buffer[4]<<10)+(in_buffer[4]<<11))-(0+(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<6)-(in_buffer[5]<<8)+(in_buffer[5]<<12))+(0-(in_buffer[6]<<1)+(in_buffer[6]<<4)-(in_buffer[6]<<6)+(in_buffer[6]<<8)+(in_buffer[6]<<9)+(in_buffer[6]<<12))+(0+(in_buffer[7]<<0)-(in_buffer[7]<<3)+(in_buffer[7]<<7)+(in_buffer[7]<<9)+(in_buffer[7]<<11)+(in_buffer[7]<<13))-(0+(in_buffer[8]<<0)-(in_buffer[8]<<2)+(in_buffer[8]<<6)-(in_buffer[8]<<8)+(in_buffer[8]<<12))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<1)+(in_buffer[9]<<6)+(in_buffer[9]<<9)+(in_buffer[9]<<11)+(in_buffer[9]<<12))-(0+(in_buffer[10]<<2)+(in_buffer[10]<<3)+(in_buffer[10]<<6)+(in_buffer[10]<<8))-(0+(in_buffer[11]<<0)+(in_buffer[11]<<2)-(in_buffer[11]<<5)-(in_buffer[11]<<8)+(in_buffer[11]<<10)+(in_buffer[11]<<11)+(in_buffer[11]<<14))-(0+(in_buffer[12]<<3)+(in_buffer[12]<<4)-(in_buffer[12]<<10)+(in_buffer[12]<<12)+(in_buffer[12]<<13))-(0-(in_buffer[13]<<0)+(in_buffer[13]<<6)+(in_buffer[13]<<7)+(in_buffer[13]<<13))-(0+(in_buffer[14]<<0)-(in_buffer[14]<<3)+(in_buffer[14]<<8))-(0+(in_buffer[15]<<5)+(in_buffer[15]<<6)+(in_buffer[15]<<9)+(in_buffer[15]<<11))+(0+(in_buffer[16]<<3)-(in_buffer[16]<<6)+(in_buffer[16]<<11))+(0+(in_buffer[17]<<3)+(in_buffer[17]<<5)+(in_buffer[17]<<9)+(in_buffer[17]<<12))+(0+(in_buffer[18]<<2)+(in_buffer[18]<<3)-(in_buffer[18]<<9)+(in_buffer[18]<<11)+(in_buffer[18]<<12))-(0-(in_buffer[19]<<0)-(in_buffer[19]<<2)-(in_buffer[19]<<4)+(in_buffer[19]<<8)+(in_buffer[19]<<9))-(0+(in_buffer[20]<<1)+(in_buffer[20]<<3)+(in_buffer[20]<<7)+(in_buffer[20]<<10))+(0+(in_buffer[21]<<1)+(in_buffer[21]<<2)+(in_buffer[21]<<5)+(in_buffer[21]<<7))+(0+(in_buffer[22]<<0)+(in_buffer[22]<<2)-(in_buffer[22]<<4)-(in_buffer[22]<<7)+(in_buffer[22]<<11))+(0+(in_buffer[23]<<0)+(in_buffer[23]<<6)+(in_buffer[23]<<7)+(in_buffer[23]<<11))-(0+(in_buffer[24]<<2)+(in_buffer[24]<<3)-(in_buffer[24]<<9)+(in_buffer[24]<<11)+(in_buffer[24]<<12))+(0-(in_buffer[25]<<0)+(in_buffer[25]<<4)+(in_buffer[25]<<5)+(in_buffer[25]<<8)+(in_buffer[25]<<12))+(0-(in_buffer[26]<<1)-(in_buffer[26]<<3)-(in_buffer[26]<<5)+(in_buffer[26]<<9)+(in_buffer[26]<<10))+(0-(in_buffer[27]<<0)-(in_buffer[27]<<2)-(in_buffer[27]<<4)+(in_buffer[27]<<8)+(in_buffer[27]<<9))+(0+(in_buffer[28]<<0)-(in_buffer[28]<<2)-(in_buffer[28]<<4)+(in_buffer[28]<<7)+(in_buffer[28]<<10)+(in_buffer[28]<<12))+(0-(in_buffer[29]<<1)+(in_buffer[29]<<11)+(in_buffer[29]<<12))-(0+(in_buffer[30]<<0)+(in_buffer[30]<<1)-(in_buffer[30]<<4)-(in_buffer[30]<<6)-(in_buffer[30]<<8)+(in_buffer[30]<<10)+(in_buffer[30]<<11))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<5)+(in_buffer[31]<<8)+(in_buffer[31]<<9)+(in_buffer[31]<<12))+(0+(in_buffer[32]<<0)+(in_buffer[32]<<6)+(in_buffer[32]<<7)+(in_buffer[32]<<11))+(0+(in_buffer[33]<<1)+(in_buffer[33]<<7)+(in_buffer[33]<<8)+(in_buffer[33]<<12))+(0+(in_buffer[34]<<1)-(in_buffer[34]<<5)-(in_buffer[34]<<10)+(in_buffer[34]<<13))+(0-(in_buffer[35]<<0)+(in_buffer[35]<<3)-(in_buffer[35]<<5)+(in_buffer[35]<<7)+(in_buffer[35]<<8)+(in_buffer[35]<<11))+(0+(in_buffer[36]<<2)+(in_buffer[36]<<4)+(in_buffer[36]<<8)+(in_buffer[36]<<11))+(0+(in_buffer[37]<<0)+(in_buffer[37]<<3)+(in_buffer[37]<<5)+(in_buffer[37]<<9)+(in_buffer[37]<<10))+(0-(in_buffer[38]<<0)+(in_buffer[38]<<5)+(in_buffer[38]<<7)+(in_buffer[38]<<8))-(0+(in_buffer[39]<<3)+(in_buffer[39]<<4)-(in_buffer[39]<<10)+(in_buffer[39]<<12)+(in_buffer[39]<<13))-(0+(in_buffer[40]<<4)-(in_buffer[40]<<7)+(in_buffer[40]<<12))+(0+(in_buffer[41]<<2)-(in_buffer[41]<<4)-(in_buffer[41]<<7)+(in_buffer[41]<<10)+(in_buffer[41]<<12))-(0+(in_buffer[42]<<3)-(in_buffer[42]<<6)+(in_buffer[42]<<11))+(0-(in_buffer[43]<<0)+(in_buffer[43]<<5)+(in_buffer[43]<<7)+(in_buffer[43]<<8))-(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<7)+(in_buffer[44]<<9)+(in_buffer[44]<<12))+(0-(in_buffer[45]<<2)-(in_buffer[45]<<4)-(in_buffer[45]<<6)+(in_buffer[45]<<10)+(in_buffer[45]<<11))+(0-(in_buffer[46]<<4)+(in_buffer[46]<<9)+(in_buffer[46]<<11)+(in_buffer[46]<<12))+(0+(in_buffer[47]<<2)+(in_buffer[47]<<4)+(in_buffer[47]<<8)+(in_buffer[47]<<11))+(0+(in_buffer[48]<<0)+(in_buffer[48]<<1)-(in_buffer[48]<<4)-(in_buffer[48]<<6)-(in_buffer[48]<<8)+(in_buffer[48]<<10)+(in_buffer[48]<<11))+(0-(in_buffer[49]<<1)+(in_buffer[49]<<4)-(in_buffer[49]<<6)+(in_buffer[49]<<8)+(in_buffer[49]<<9)+(in_buffer[49]<<12))-(0+(in_buffer[50]<<3)-(in_buffer[50]<<6)+(in_buffer[50]<<11))-(0+(in_buffer[51]<<6)+(in_buffer[51]<<7)+(in_buffer[51]<<10)+(in_buffer[51]<<12))+(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)-(in_buffer[52]<<4)-(in_buffer[52]<<6)+(in_buffer[52]<<11)+(in_buffer[52]<<12))+(0-(in_buffer[53]<<0)-(in_buffer[53]<<2)+(in_buffer[53]<<5)+(in_buffer[53]<<11))-(0+(in_buffer[54]<<1)+(in_buffer[54]<<2)-(in_buffer[54]<<6)+(in_buffer[54]<<13))+(0+(in_buffer[55]<<0)-(in_buffer[55]<<2)-(in_buffer[55]<<5)+(in_buffer[55]<<8)+(in_buffer[55]<<10))-(0+(in_buffer[56]<<1)+(in_buffer[56]<<5)-(in_buffer[56]<<8)+(in_buffer[56]<<11))-(0+(in_buffer[57]<<3)+(in_buffer[57]<<4)+(in_buffer[57]<<7)+(in_buffer[57]<<9))-(0-(in_buffer[58]<<1)+(in_buffer[58]<<5)+(in_buffer[58]<<6)+(in_buffer[58]<<9)+(in_buffer[58]<<13))-(0+(in_buffer[59]<<1)+(in_buffer[59]<<3)-(in_buffer[59]<<5)-(in_buffer[59]<<8)+(in_buffer[59]<<12))+(0-(in_buffer[60]<<2)-(in_buffer[60]<<5)+(in_buffer[60]<<8)+(in_buffer[60]<<12))+(0+(in_buffer[61]<<1)+(in_buffer[61]<<4)+(in_buffer[61]<<8)+(in_buffer[61]<<13))-(0+(in_buffer[62]<<1)+(in_buffer[62]<<2)+(in_buffer[62]<<5)+(in_buffer[62]<<7))-(0+(in_buffer[63]<<0)-(in_buffer[63]<<3)+(in_buffer[63]<<8))-(0+(in_buffer[64]<<0)+(in_buffer[64]<<1)-(in_buffer[64]<<4)-(in_buffer[64]<<6)-(in_buffer[64]<<8)+(in_buffer[64]<<10)+(in_buffer[64]<<11))-(0+(in_buffer[65]<<2)+(in_buffer[65]<<6)-(in_buffer[65]<<9)+(in_buffer[65]<<12))+(0+(in_buffer[66]<<1)+(in_buffer[66]<<3)-(in_buffer[66]<<5)-(in_buffer[66]<<8)+(in_buffer[66]<<12))+(0+(in_buffer[67]<<1)+(in_buffer[67]<<7)+(in_buffer[67]<<8)+(in_buffer[67]<<12))-(0+(in_buffer[68]<<0)+(in_buffer[68]<<2)+(in_buffer[68]<<6)+(in_buffer[68]<<9))+(0+(in_buffer[69]<<1)-(in_buffer[69]<<4)+(in_buffer[69]<<9))-(0+(in_buffer[70]<<0)+(in_buffer[70]<<4)-(in_buffer[70]<<7)+(in_buffer[70]<<10))+(0-(in_buffer[71]<<0)+(in_buffer[71]<<4)-(in_buffer[71]<<6)-(in_buffer[71]<<8)+(in_buffer[71]<<11))+(0-(in_buffer[72]<<0)+(in_buffer[72]<<4)-(in_buffer[72]<<6)-(in_buffer[72]<<8)+(in_buffer[72]<<11))+(0-(in_buffer[73]<<1)+(in_buffer[73]<<4)-(in_buffer[73]<<6)+(in_buffer[73]<<8)+(in_buffer[73]<<9)+(in_buffer[73]<<12))-(0+(in_buffer[74]<<0)+(in_buffer[74]<<6)+(in_buffer[74]<<7)+(in_buffer[74]<<11))-(0+(in_buffer[75]<<5)+(in_buffer[75]<<6)+(in_buffer[75]<<9)+(in_buffer[75]<<11))+(0+(in_buffer[76]<<1)-(in_buffer[76]<<3)+(in_buffer[76]<<7)-(in_buffer[76]<<9)+(in_buffer[76]<<13))-(0+(in_buffer[77]<<1)+(in_buffer[77]<<3)+(in_buffer[77]<<7)+(in_buffer[77]<<10))-(0+(in_buffer[78]<<2)-(in_buffer[78]<<5)+(in_buffer[78]<<10))-(0-(in_buffer[79]<<0)+(in_buffer[79]<<3)-(in_buffer[79]<<6)+(in_buffer[79]<<10)+(in_buffer[79]<<12))+(0+(in_buffer[80]<<0)+(in_buffer[80]<<1)-(in_buffer[80]<<7)+(in_buffer[80]<<9)+(in_buffer[80]<<10))-(0+(in_buffer[81]<<2)+(in_buffer[81]<<3)+(in_buffer[81]<<6)+(in_buffer[81]<<8))-(0+(in_buffer[82]<<1)+(in_buffer[82]<<5)-(in_buffer[82]<<8)+(in_buffer[82]<<11))-(0-(in_buffer[83]<<0)+(in_buffer[83]<<3)-(in_buffer[83]<<5)+(in_buffer[83]<<7)+(in_buffer[83]<<8)+(in_buffer[83]<<11))+(0+(in_buffer[84]<<1)+(in_buffer[84]<<2)+(in_buffer[84]<<5)+(in_buffer[84]<<7))-(0+(in_buffer[85]<<0)+(in_buffer[85]<<2)+(in_buffer[85]<<3)+(in_buffer[85]<<9)+(in_buffer[85]<<11))+(0-(in_buffer[86]<<0)-(in_buffer[86]<<3)+(in_buffer[86]<<6)+(in_buffer[86]<<10))-(0+(in_buffer[87]<<0)-(in_buffer[87]<<3)+(in_buffer[87]<<8))+(0+(in_buffer[88]<<2)+(in_buffer[88]<<3)+(in_buffer[88]<<6)+(in_buffer[88]<<8))-(0-(in_buffer[89]<<0)+(in_buffer[89]<<2)+(in_buffer[89]<<3)+(in_buffer[89]<<6)+(in_buffer[89]<<8)+(in_buffer[89]<<10)+(in_buffer[89]<<11))-(0-(in_buffer[90]<<0)-(in_buffer[90]<<2)-(in_buffer[90]<<4)-(in_buffer[90]<<6)+(in_buffer[90]<<11)+(in_buffer[90]<<12))+(0-(in_buffer[91]<<0)+(in_buffer[91]<<3)+(in_buffer[91]<<4)+(in_buffer[91]<<7)-(in_buffer[91]<<9)+(in_buffer[91]<<12))+(0-(in_buffer[92]<<1)+(in_buffer[92]<<6)+(in_buffer[92]<<8)+(in_buffer[92]<<9))-(0+(in_buffer[93]<<0)+(in_buffer[93]<<1)+(in_buffer[93]<<4)+(in_buffer[93]<<6))-(0-(in_buffer[94]<<2)+(in_buffer[94]<<7)+(in_buffer[94]<<9)+(in_buffer[94]<<10))-(0+(in_buffer[95]<<1)+(in_buffer[95]<<2)-(in_buffer[95]<<8)+(in_buffer[95]<<10)+(in_buffer[95]<<11))-(0-(in_buffer[96]<<0)+(in_buffer[96]<<6)+(in_buffer[96]<<7)+(in_buffer[96]<<13))-(0+(in_buffer[97]<<0)+(in_buffer[97]<<4)+(in_buffer[97]<<6)+(in_buffer[97]<<11)+(in_buffer[97]<<12))+(0+(in_buffer[98]<<2)-(in_buffer[98]<<5)+(in_buffer[98]<<10))-(0+(in_buffer[99]<<0)-(in_buffer[99]<<2)+(in_buffer[99]<<6)-(in_buffer[99]<<8)+(in_buffer[99]<<12))-(0+(in_buffer[100]<<0)-(in_buffer[100]<<2)-(in_buffer[100]<<4)+(in_buffer[100]<<7)+(in_buffer[100]<<10)+(in_buffer[100]<<12))-(0-(in_buffer[101]<<0)+(in_buffer[101]<<3)-(in_buffer[101]<<6)+(in_buffer[101]<<10)+(in_buffer[101]<<12))+(0+(in_buffer[102]<<0)+(in_buffer[102]<<2)+(in_buffer[102]<<3)-(in_buffer[102]<<6)-(in_buffer[102]<<8)+(in_buffer[102]<<13))+(0+(in_buffer[103]<<0)+(in_buffer[103]<<2)+(in_buffer[103]<<3)-(in_buffer[103]<<6)-(in_buffer[103]<<8)+(in_buffer[103]<<13))+(0-(in_buffer[104]<<0)+(in_buffer[104]<<5)+(in_buffer[104]<<6)-(in_buffer[104]<<9)+(in_buffer[104]<<11)+(in_buffer[104]<<12))-(0+(in_buffer[105]<<2)-(in_buffer[105]<<5)+(in_buffer[105]<<10))+(0-(in_buffer[106]<<1)+(in_buffer[106]<<6)+(in_buffer[106]<<8)+(in_buffer[106]<<9))-(0+(in_buffer[107]<<0)-(in_buffer[107]<<4)-(in_buffer[107]<<9)+(in_buffer[107]<<12))-(0+(in_buffer[108]<<0)-(in_buffer[108]<<3)-(in_buffer[108]<<6)-(in_buffer[108]<<9)+(in_buffer[108]<<11)+(in_buffer[108]<<12))+(0+(in_buffer[109]<<0)+(in_buffer[109]<<1)-(in_buffer[109]<<4)-(in_buffer[109]<<7)+(in_buffer[109]<<13))+(0+(in_buffer[110]<<0)+(in_buffer[110]<<3)+(in_buffer[110]<<5)+(in_buffer[110]<<9)+(in_buffer[110]<<10))-(0-(in_buffer[111]<<0)-(in_buffer[111]<<2)+(in_buffer[111]<<7)+(in_buffer[111]<<9)+(in_buffer[111]<<12))-(0-(in_buffer[112]<<1)+(in_buffer[112]<<5)-(in_buffer[112]<<7)-(in_buffer[112]<<9)+(in_buffer[112]<<12))+(0+(in_buffer[113]<<3)+(in_buffer[113]<<7)-(in_buffer[113]<<10)+(in_buffer[113]<<13))+(0+(in_buffer[114]<<0)-(in_buffer[114]<<3)-(in_buffer[114]<<5)-(in_buffer[114]<<7)+(in_buffer[114]<<10)+(in_buffer[114]<<11))+(0+(in_buffer[115]<<0)-(in_buffer[115]<<2)-(in_buffer[115]<<5)+(in_buffer[115]<<8)+(in_buffer[115]<<10))-(0-(in_buffer[116]<<0)+(in_buffer[116]<<3)+(in_buffer[116]<<4)+(in_buffer[116]<<7)-(in_buffer[116]<<9)+(in_buffer[116]<<12))+(0+(in_buffer[117]<<0)+(in_buffer[117]<<2)+(in_buffer[117]<<4)-(in_buffer[117]<<6)+(in_buffer[117]<<9)+(in_buffer[117]<<12))+(0-(in_buffer[118]<<3)-(in_buffer[118]<<5)-(in_buffer[118]<<7)+(in_buffer[118]<<11)+(in_buffer[118]<<12))-(0-(in_buffer[119]<<1)+(in_buffer[119]<<4)-(in_buffer[119]<<6)+(in_buffer[119]<<8)+(in_buffer[119]<<9)+(in_buffer[119]<<12))-(0+(in_buffer[120]<<0)-(in_buffer[120]<<2)-(in_buffer[120]<<5)+(in_buffer[120]<<8)+(in_buffer[120]<<10));
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
wire signed [DATA_WIDTH-1:0]   weight_bias10;
wire signed [DATA_WIDTH-1:0]   weight_bias11;
wire signed [DATA_WIDTH-1:0]   weight_bias12;
wire signed [DATA_WIDTH-1:0]   weight_bias13;
wire signed [DATA_WIDTH-1:0]   weight_bias14;
wire signed [DATA_WIDTH-1:0]   weight_bias15;
wire signed [DATA_WIDTH-1:0]   weight_bias16;
wire signed [DATA_WIDTH-1:0]   weight_bias17;
wire signed [DATA_WIDTH-1:0]   weight_bias18;
wire signed [DATA_WIDTH-1:0]   weight_bias19;
wire signed [DATA_WIDTH-1:0]   weight_bias20;
wire signed [DATA_WIDTH-1:0]   weight_bias21;
wire signed [DATA_WIDTH-1:0]   weight_bias22;
wire signed [DATA_WIDTH-1:0]   weight_bias23;
wire signed [DATA_WIDTH-1:0]   weight_bias24;
wire signed [DATA_WIDTH-1:0]   weight_bias25;
wire signed [DATA_WIDTH-1:0]   weight_bias26;
wire signed [DATA_WIDTH-1:0]   weight_bias27;
wire signed [DATA_WIDTH-1:0]   weight_bias28;
wire signed [DATA_WIDTH-1:0]   weight_bias29;
wire signed [DATA_WIDTH-1:0]   weight_bias30;
wire signed [DATA_WIDTH-1:0]   weight_bias31;
assign weight_bias0=in_buffer_weight0+(1577);
assign weight_bias1=in_buffer_weight1+(4980);
assign weight_bias2=in_buffer_weight2+(-5727);
assign weight_bias3=in_buffer_weight3+(7221);
assign weight_bias4=in_buffer_weight4+(-1494);
assign weight_bias5=in_buffer_weight5+(-6889);
assign weight_bias6=in_buffer_weight6+(6889);
assign weight_bias7=in_buffer_weight7+(6142);
assign weight_bias8=in_buffer_weight8+(-1411);
assign weight_bias9=in_buffer_weight9+(0);
assign weight_bias10=in_buffer_weight10+(2739);
assign weight_bias11=in_buffer_weight11+(-913);
assign weight_bias12=in_buffer_weight12+(7636);
assign weight_bias13=in_buffer_weight13+(-1577);
assign weight_bias14=in_buffer_weight14+(3237);
assign weight_bias15=in_buffer_weight15+(-5810);
assign weight_bias16=in_buffer_weight16+(-581);
assign weight_bias17=in_buffer_weight17+(-2739);
assign weight_bias18=in_buffer_weight18+(-166);
assign weight_bias19=in_buffer_weight19+(7636);
assign weight_bias20=in_buffer_weight20+(2905);
assign weight_bias21=in_buffer_weight21+(2158);
assign weight_bias22=in_buffer_weight22+(-581);
assign weight_bias23=in_buffer_weight23+(-747);
assign weight_bias24=in_buffer_weight24+(5063);
assign weight_bias25=in_buffer_weight25+(8300);
assign weight_bias26=in_buffer_weight26+(-2241);
assign weight_bias27=in_buffer_weight27+(-913);
assign weight_bias28=in_buffer_weight28+(1826);
assign weight_bias29=in_buffer_weight29+(3403);
assign weight_bias30=in_buffer_weight30+(10209);
assign weight_bias31=in_buffer_weight31+(996);
wire signed [DATA_WIDTH-1:0]   bias_relu0;
wire signed [DATA_WIDTH-1:0]   bias_relu1;
wire signed [DATA_WIDTH-1:0]   bias_relu2;
wire signed [DATA_WIDTH-1:0]   bias_relu3;
wire signed [DATA_WIDTH-1:0]   bias_relu4;
wire signed [DATA_WIDTH-1:0]   bias_relu5;
wire signed [DATA_WIDTH-1:0]   bias_relu6;
wire signed [DATA_WIDTH-1:0]   bias_relu7;
wire signed [DATA_WIDTH-1:0]   bias_relu8;
wire signed [DATA_WIDTH-1:0]   bias_relu9;
wire signed [DATA_WIDTH-1:0]   bias_relu10;
wire signed [DATA_WIDTH-1:0]   bias_relu11;
wire signed [DATA_WIDTH-1:0]   bias_relu12;
wire signed [DATA_WIDTH-1:0]   bias_relu13;
wire signed [DATA_WIDTH-1:0]   bias_relu14;
wire signed [DATA_WIDTH-1:0]   bias_relu15;
wire signed [DATA_WIDTH-1:0]   bias_relu16;
wire signed [DATA_WIDTH-1:0]   bias_relu17;
wire signed [DATA_WIDTH-1:0]   bias_relu18;
wire signed [DATA_WIDTH-1:0]   bias_relu19;
wire signed [DATA_WIDTH-1:0]   bias_relu20;
wire signed [DATA_WIDTH-1:0]   bias_relu21;
wire signed [DATA_WIDTH-1:0]   bias_relu22;
wire signed [DATA_WIDTH-1:0]   bias_relu23;
wire signed [DATA_WIDTH-1:0]   bias_relu24;
wire signed [DATA_WIDTH-1:0]   bias_relu25;
wire signed [DATA_WIDTH-1:0]   bias_relu26;
wire signed [DATA_WIDTH-1:0]   bias_relu27;
wire signed [DATA_WIDTH-1:0]   bias_relu28;
wire signed [DATA_WIDTH-1:0]   bias_relu29;
wire signed [DATA_WIDTH-1:0]   bias_relu30;
wire signed [DATA_WIDTH-1:0]   bias_relu31;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign layer_out={bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule