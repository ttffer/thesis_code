module an_decorder_n13_testbench ();
	
	
	an_decoder_n13

endmodule